module VTASim(
  input   clock,
  input   reset,
  output  sim_wait
);
  wire  sim_clock; // @[SimShell.scala 55:19]
  wire  sim_reset; // @[SimShell.scala 55:19]
  wire  sim_dpi_wait; // @[SimShell.scala 55:19]
  VTASimDPI sim ( // @[SimShell.scala 55:19]
    .clock(sim_clock),
    .reset(sim_reset),
    .dpi_wait(sim_dpi_wait)
  );
  assign sim_wait = sim_dpi_wait; // @[SimShell.scala 58:12]
  assign sim_clock = clock; // @[SimShell.scala 57:16]
  assign sim_reset = reset; // @[SimShell.scala 56:16]
endmodule
module VTAHostDPIToAXI(
  input         clock,
  input         reset,
  input         io_dpi_req_valid,
  input         io_dpi_req_opcode,
  input  [31:0] io_dpi_req_addr,
  input  [31:0] io_dpi_req_value,
  output        io_dpi_req_deq,
  output        io_dpi_resp_valid,
  output [31:0] io_dpi_resp_bits,
  input         io_axi_aw_ready,
  output        io_axi_aw_valid,
  output [31:0] io_axi_aw_bits_addr,
  input         io_axi_w_ready,
  output        io_axi_w_valid,
  output [63:0] io_axi_w_bits_data,
  output        io_axi_b_ready,
  input         io_axi_b_valid,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [31:0] io_axi_ar_bits_addr,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [63:0] io_axi_r_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] addr; // @[VTAHostDPI.scala 69:21]
  reg [31:0] data; // @[VTAHostDPI.scala 70:21]
  reg [2:0] state; // @[VTAHostDPI.scala 73:22]
  wire  _T_2 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_6 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_8 = state == 3'h0; // @[VTAHostDPI.scala 112:14]
  wire  _T_9 = _T_8 & io_dpi_req_valid; // @[VTAHostDPI.scala 112:24]
  wire  _T_10 = state == 3'h3; // @[VTAHostDPI.scala 117:28]
  wire  _T_13 = state == 3'h1; // @[VTAHostDPI.scala 124:28]
  wire  _T_16 = _T_13 & io_axi_ar_ready; // @[VTAHostDPI.scala 128:45]
  wire  _T_18 = _T_10 & io_axi_aw_ready; // @[VTAHostDPI.scala 128:91]
  assign io_dpi_req_deq = _T_16 | _T_18; // @[VTAHostDPI.scala 128:18]
  assign io_dpi_resp_valid = io_axi_r_valid; // @[VTAHostDPI.scala 129:21]
  assign io_dpi_resp_bits = io_axi_r_bits_data[31:0]; // @[VTAHostDPI.scala 130:20]
  assign io_axi_aw_valid = state == 3'h3; // @[VTAHostDPI.scala 117:19]
  assign io_axi_aw_bits_addr = addr; // @[VTAHostDPI.scala 118:23]
  assign io_axi_w_valid = state == 3'h4; // @[VTAHostDPI.scala 119:18]
  assign io_axi_w_bits_data = {{32'd0}, data}; // @[VTAHostDPI.scala 120:22]
  assign io_axi_b_ready = state == 3'h5; // @[VTAHostDPI.scala 122:18]
  assign io_axi_ar_valid = state == 3'h1; // @[VTAHostDPI.scala 124:19]
  assign io_axi_ar_bits_addr = addr; // @[VTAHostDPI.scala 125:23]
  assign io_axi_r_ready = state == 3'h2; // @[VTAHostDPI.scala 126:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  data = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr <= 32'h0;
    end else if (_T_9) begin
      addr <= io_dpi_req_addr;
    end
    if (reset) begin
      data <= 32'h0;
    end else if (_T_9) begin
      data <= io_dpi_req_value;
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_2) begin
      if (io_dpi_req_valid) begin
        if (io_dpi_req_opcode) begin
          state <= 3'h3;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (_T_3) begin
      if (io_axi_ar_ready) begin
        state <= 3'h2;
      end
    end else if (_T_4) begin
      if (io_axi_r_valid) begin
        state <= 3'h0;
      end
    end else if (_T_5) begin
      if (io_axi_aw_ready) begin
        state <= 3'h4;
      end
    end else if (_T_6) begin
      if (io_axi_w_ready) begin
        state <= 3'h5;
      end
    end else if (_T_7) begin
      if (io_axi_b_valid) begin
        state <= 3'h0;
      end
    end
  end
endmodule
module VTAHost(
  input         clock,
  input         reset,
  input         io_axi_aw_ready,
  output        io_axi_aw_valid,
  output [31:0] io_axi_aw_bits_addr,
  input         io_axi_w_ready,
  output        io_axi_w_valid,
  output [63:0] io_axi_w_bits_data,
  output        io_axi_b_ready,
  input         io_axi_b_valid,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [31:0] io_axi_ar_bits_addr,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [63:0] io_axi_r_bits_data
);
  wire  host_dpi_clock; // @[SimShell.scala 20:24]
  wire  host_dpi_reset; // @[SimShell.scala 20:24]
  wire  host_dpi_dpi_req_valid; // @[SimShell.scala 20:24]
  wire  host_dpi_dpi_req_opcode; // @[SimShell.scala 20:24]
  wire [31:0] host_dpi_dpi_req_addr; // @[SimShell.scala 20:24]
  wire [31:0] host_dpi_dpi_req_value; // @[SimShell.scala 20:24]
  wire  host_dpi_dpi_req_deq; // @[SimShell.scala 20:24]
  wire  host_dpi_dpi_resp_valid; // @[SimShell.scala 20:24]
  wire [31:0] host_dpi_dpi_resp_bits; // @[SimShell.scala 20:24]
  wire  host_axi_clock; // @[SimShell.scala 21:24]
  wire  host_axi_reset; // @[SimShell.scala 21:24]
  wire  host_axi_io_dpi_req_valid; // @[SimShell.scala 21:24]
  wire  host_axi_io_dpi_req_opcode; // @[SimShell.scala 21:24]
  wire [31:0] host_axi_io_dpi_req_addr; // @[SimShell.scala 21:24]
  wire [31:0] host_axi_io_dpi_req_value; // @[SimShell.scala 21:24]
  wire  host_axi_io_dpi_req_deq; // @[SimShell.scala 21:24]
  wire  host_axi_io_dpi_resp_valid; // @[SimShell.scala 21:24]
  wire [31:0] host_axi_io_dpi_resp_bits; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_aw_ready; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_aw_valid; // @[SimShell.scala 21:24]
  wire [31:0] host_axi_io_axi_aw_bits_addr; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_w_ready; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_w_valid; // @[SimShell.scala 21:24]
  wire [63:0] host_axi_io_axi_w_bits_data; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_b_ready; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_b_valid; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_ar_ready; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_ar_valid; // @[SimShell.scala 21:24]
  wire [31:0] host_axi_io_axi_ar_bits_addr; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_r_ready; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_r_valid; // @[SimShell.scala 21:24]
  wire [63:0] host_axi_io_axi_r_bits_data; // @[SimShell.scala 21:24]
  VTAHostDPI host_dpi ( // @[SimShell.scala 20:24]
    .clock(host_dpi_clock),
    .reset(host_dpi_reset),
    .dpi_req_valid(host_dpi_dpi_req_valid),
    .dpi_req_opcode(host_dpi_dpi_req_opcode),
    .dpi_req_addr(host_dpi_dpi_req_addr),
    .dpi_req_value(host_dpi_dpi_req_value),
    .dpi_req_deq(host_dpi_dpi_req_deq),
    .dpi_resp_valid(host_dpi_dpi_resp_valid),
    .dpi_resp_bits(host_dpi_dpi_resp_bits)
  );
  VTAHostDPIToAXI host_axi ( // @[SimShell.scala 21:24]
    .clock(host_axi_clock),
    .reset(host_axi_reset),
    .io_dpi_req_valid(host_axi_io_dpi_req_valid),
    .io_dpi_req_opcode(host_axi_io_dpi_req_opcode),
    .io_dpi_req_addr(host_axi_io_dpi_req_addr),
    .io_dpi_req_value(host_axi_io_dpi_req_value),
    .io_dpi_req_deq(host_axi_io_dpi_req_deq),
    .io_dpi_resp_valid(host_axi_io_dpi_resp_valid),
    .io_dpi_resp_bits(host_axi_io_dpi_resp_bits),
    .io_axi_aw_ready(host_axi_io_axi_aw_ready),
    .io_axi_aw_valid(host_axi_io_axi_aw_valid),
    .io_axi_aw_bits_addr(host_axi_io_axi_aw_bits_addr),
    .io_axi_w_ready(host_axi_io_axi_w_ready),
    .io_axi_w_valid(host_axi_io_axi_w_valid),
    .io_axi_w_bits_data(host_axi_io_axi_w_bits_data),
    .io_axi_b_ready(host_axi_io_axi_b_ready),
    .io_axi_b_valid(host_axi_io_axi_b_valid),
    .io_axi_ar_ready(host_axi_io_axi_ar_ready),
    .io_axi_ar_valid(host_axi_io_axi_ar_valid),
    .io_axi_ar_bits_addr(host_axi_io_axi_ar_bits_addr),
    .io_axi_r_ready(host_axi_io_axi_r_ready),
    .io_axi_r_valid(host_axi_io_axi_r_valid),
    .io_axi_r_bits_data(host_axi_io_axi_r_bits_data)
  );
  assign io_axi_aw_valid = host_axi_io_axi_aw_valid; // @[SimShell.scala 25:10]
  assign io_axi_aw_bits_addr = host_axi_io_axi_aw_bits_addr; // @[SimShell.scala 25:10]
  assign io_axi_w_valid = host_axi_io_axi_w_valid; // @[SimShell.scala 25:10]
  assign io_axi_w_bits_data = host_axi_io_axi_w_bits_data; // @[SimShell.scala 25:10]
  assign io_axi_b_ready = host_axi_io_axi_b_ready; // @[SimShell.scala 25:10]
  assign io_axi_ar_valid = host_axi_io_axi_ar_valid; // @[SimShell.scala 25:10]
  assign io_axi_ar_bits_addr = host_axi_io_axi_ar_bits_addr; // @[SimShell.scala 25:10]
  assign io_axi_r_ready = host_axi_io_axi_r_ready; // @[SimShell.scala 25:10]
  assign host_dpi_clock = clock; // @[SimShell.scala 23:21]
  assign host_dpi_reset = reset; // @[SimShell.scala 22:21]
  assign host_dpi_dpi_req_deq = host_axi_io_dpi_req_deq; // @[SimShell.scala 24:19]
  assign host_dpi_dpi_resp_valid = host_axi_io_dpi_resp_valid; // @[SimShell.scala 24:19]
  assign host_dpi_dpi_resp_bits = host_axi_io_dpi_resp_bits; // @[SimShell.scala 24:19]
  assign host_axi_clock = clock;
  assign host_axi_reset = reset;
  assign host_axi_io_dpi_req_valid = host_dpi_dpi_req_valid; // @[SimShell.scala 24:19]
  assign host_axi_io_dpi_req_opcode = host_dpi_dpi_req_opcode; // @[SimShell.scala 24:19]
  assign host_axi_io_dpi_req_addr = host_dpi_dpi_req_addr; // @[SimShell.scala 24:19]
  assign host_axi_io_dpi_req_value = host_dpi_dpi_req_value; // @[SimShell.scala 24:19]
  assign host_axi_io_axi_aw_ready = io_axi_aw_ready; // @[SimShell.scala 25:10]
  assign host_axi_io_axi_w_ready = io_axi_w_ready; // @[SimShell.scala 25:10]
  assign host_axi_io_axi_b_valid = io_axi_b_valid; // @[SimShell.scala 25:10]
  assign host_axi_io_axi_ar_ready = io_axi_ar_ready; // @[SimShell.scala 25:10]
  assign host_axi_io_axi_r_valid = io_axi_r_valid; // @[SimShell.scala 25:10]
  assign host_axi_io_axi_r_bits_data = io_axi_r_bits_data; // @[SimShell.scala 25:10]
endmodule
module VTAMemDPIToAXI(
  input         clock,
  input         reset,
  output        io_dpi_req_valid,
  output        io_dpi_req_opcode,
  output [31:0] io_dpi_req_len,
  output [63:0] io_dpi_req_addr,
  output        io_dpi_wr_valid,
  output [63:0] io_dpi_wr_bits,
  output        io_dpi_rd_ready,
  input         io_dpi_rd_valid,
  input  [63:0] io_dpi_rd_bits,
  output        io_axi_aw_ready,
  input         io_axi_aw_valid,
  input  [31:0] io_axi_aw_bits_addr,
  input  [31:0] io_axi_aw_bits_len,
  output        io_axi_w_ready,
  input         io_axi_w_valid,
  input  [63:0] io_axi_w_bits_data,
  input         io_axi_w_bits_last,
  input         io_axi_b_ready,
  output        io_axi_b_valid,
  output        io_axi_ar_ready,
  input         io_axi_ar_valid,
  input  [31:0] io_axi_ar_bits_addr,
  input  [31:0] io_axi_ar_bits_len,
  input         io_axi_r_ready,
  output        io_axi_r_valid,
  output [63:0] io_axi_r_bits_data,
  output        io_axi_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  opcode; // @[VTAMemDPI.scala 85:23]
  reg [31:0] len; // @[VTAMemDPI.scala 86:20]
  reg [63:0] addr; // @[VTAMemDPI.scala 87:21]
  reg [2:0] state; // @[VTAMemDPI.scala 90:22]
  wire  _T_2 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = io_axi_r_ready & io_dpi_rd_valid; // @[VTAMemDPI.scala 106:27]
  wire  _T_6 = len == 32'h0; // @[VTAMemDPI.scala 106:53]
  wire  _T_7 = _T_5 & _T_6; // @[VTAMemDPI.scala 106:46]
  wire  _T_8 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_10 = io_axi_w_valid & io_axi_w_bits_last; // @[VTAMemDPI.scala 116:27]
  wire  _T_11 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = state == 3'h0; // @[VTAMemDPI.scala 127:14]
  wire  _GEN_13 = io_axi_aw_valid | opcode; // @[VTAMemDPI.scala 132:33]
  wire  _T_13 = state == 3'h2; // @[VTAMemDPI.scala 138:20]
  wire  _T_15 = len != 32'h0; // @[VTAMemDPI.scala 139:51]
  wire  _T_16 = _T_5 & _T_15; // @[VTAMemDPI.scala 139:44]
  wire [31:0] _T_18 = len - 32'h1; // @[VTAMemDPI.scala 140:18]
  wire  _T_19 = state == 3'h1; // @[VTAMemDPI.scala 144:30]
  wire  _T_20 = _T_19 & io_axi_ar_valid; // @[VTAMemDPI.scala 144:47]
  wire  _T_21 = state == 3'h3; // @[VTAMemDPI.scala 144:75]
  wire  _T_22 = _T_21 & io_axi_aw_valid; // @[VTAMemDPI.scala 144:93]
  wire  _T_31 = state == 3'h4; // @[VTAMemDPI.scala 160:28]
  assign io_dpi_req_valid = _T_20 | _T_22; // @[VTAMemDPI.scala 144:20]
  assign io_dpi_req_opcode = opcode; // @[VTAMemDPI.scala 145:21]
  assign io_dpi_req_len = len; // @[VTAMemDPI.scala 146:18]
  assign io_dpi_req_addr = addr; // @[VTAMemDPI.scala 147:19]
  assign io_dpi_wr_valid = _T_31 & io_axi_w_valid; // @[VTAMemDPI.scala 160:19]
  assign io_dpi_wr_bits = io_axi_w_bits_data; // @[VTAMemDPI.scala 161:18]
  assign io_dpi_rd_ready = _T_13 & io_axi_r_ready; // @[VTAMemDPI.scala 158:19]
  assign io_axi_aw_ready = state == 3'h3; // @[VTAMemDPI.scala 150:19]
  assign io_axi_w_ready = state == 3'h4; // @[VTAMemDPI.scala 162:18]
  assign io_axi_b_valid = state == 3'h5; // @[VTAMemDPI.scala 164:18]
  assign io_axi_ar_ready = state == 3'h1; // @[VTAMemDPI.scala 149:19]
  assign io_axi_r_valid = _T_13 & io_dpi_rd_valid; // @[VTAMemDPI.scala 152:18]
  assign io_axi_r_bits_data = io_dpi_rd_bits; // @[VTAMemDPI.scala 153:22]
  assign io_axi_r_bits_last = len == 32'h0; // @[VTAMemDPI.scala 154:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  opcode = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  len = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  addr = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      opcode <= 1'h0;
    end else if (_T_12) begin
      if (io_axi_ar_valid) begin
        opcode <= 1'h0;
      end else begin
        opcode <= _GEN_13;
      end
    end
    if (reset) begin
      len <= 32'h0;
    end else if (_T_12) begin
      if (io_axi_ar_valid) begin
        len <= io_axi_ar_bits_len;
      end else if (io_axi_aw_valid) begin
        len <= io_axi_aw_bits_len;
      end
    end else if (_T_13) begin
      if (_T_16) begin
        len <= _T_18;
      end
    end
    if (reset) begin
      addr <= 64'h0;
    end else if (_T_12) begin
      if (io_axi_ar_valid) begin
        addr <= {{32'd0}, io_axi_ar_bits_addr};
      end else if (io_axi_aw_valid) begin
        addr <= {{32'd0}, io_axi_aw_bits_addr};
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_2) begin
      if (io_axi_ar_valid) begin
        state <= 3'h1;
      end else if (io_axi_aw_valid) begin
        state <= 3'h3;
      end
    end else if (_T_3) begin
      if (io_axi_ar_valid) begin
        state <= 3'h2;
      end
    end else if (_T_4) begin
      if (_T_7) begin
        state <= 3'h0;
      end
    end else if (_T_8) begin
      if (io_axi_aw_valid) begin
        state <= 3'h4;
      end
    end else if (_T_9) begin
      if (_T_10) begin
        state <= 3'h5;
      end
    end else if (_T_11) begin
      if (io_axi_b_ready) begin
        state <= 3'h0;
      end
    end
  end
endmodule
module VTAMem(
  input         clock,
  input         reset,
  output        io_axi_aw_ready,
  input         io_axi_aw_valid,
  input  [31:0] io_axi_aw_bits_addr,
  input  [31:0] io_axi_aw_bits_len,
  output        io_axi_w_ready,
  input         io_axi_w_valid,
  input  [63:0] io_axi_w_bits_data,
  input         io_axi_w_bits_last,
  input         io_axi_b_ready,
  output        io_axi_b_valid,
  output        io_axi_ar_ready,
  input         io_axi_ar_valid,
  input  [31:0] io_axi_ar_bits_addr,
  input  [31:0] io_axi_ar_bits_len,
  input         io_axi_r_ready,
  output        io_axi_r_valid,
  output [63:0] io_axi_r_bits_data,
  output        io_axi_r_bits_last
);
  wire  mem_dpi_clock; // @[SimShell.scala 38:23]
  wire  mem_dpi_reset; // @[SimShell.scala 38:23]
  wire  mem_dpi_dpi_req_valid; // @[SimShell.scala 38:23]
  wire  mem_dpi_dpi_req_opcode; // @[SimShell.scala 38:23]
  wire [31:0] mem_dpi_dpi_req_len; // @[SimShell.scala 38:23]
  wire [63:0] mem_dpi_dpi_req_addr; // @[SimShell.scala 38:23]
  wire  mem_dpi_dpi_wr_valid; // @[SimShell.scala 38:23]
  wire [63:0] mem_dpi_dpi_wr_bits; // @[SimShell.scala 38:23]
  wire  mem_dpi_dpi_rd_ready; // @[SimShell.scala 38:23]
  wire  mem_dpi_dpi_rd_valid; // @[SimShell.scala 38:23]
  wire [63:0] mem_dpi_dpi_rd_bits; // @[SimShell.scala 38:23]
  wire  mem_axi_clock; // @[SimShell.scala 39:23]
  wire  mem_axi_reset; // @[SimShell.scala 39:23]
  wire  mem_axi_io_dpi_req_valid; // @[SimShell.scala 39:23]
  wire  mem_axi_io_dpi_req_opcode; // @[SimShell.scala 39:23]
  wire [31:0] mem_axi_io_dpi_req_len; // @[SimShell.scala 39:23]
  wire [63:0] mem_axi_io_dpi_req_addr; // @[SimShell.scala 39:23]
  wire  mem_axi_io_dpi_wr_valid; // @[SimShell.scala 39:23]
  wire [63:0] mem_axi_io_dpi_wr_bits; // @[SimShell.scala 39:23]
  wire  mem_axi_io_dpi_rd_ready; // @[SimShell.scala 39:23]
  wire  mem_axi_io_dpi_rd_valid; // @[SimShell.scala 39:23]
  wire [63:0] mem_axi_io_dpi_rd_bits; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_aw_ready; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_aw_valid; // @[SimShell.scala 39:23]
  wire [31:0] mem_axi_io_axi_aw_bits_addr; // @[SimShell.scala 39:23]
  wire [31:0] mem_axi_io_axi_aw_bits_len; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_w_ready; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_w_valid; // @[SimShell.scala 39:23]
  wire [63:0] mem_axi_io_axi_w_bits_data; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_w_bits_last; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_b_ready; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_b_valid; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_ar_ready; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_ar_valid; // @[SimShell.scala 39:23]
  wire [31:0] mem_axi_io_axi_ar_bits_addr; // @[SimShell.scala 39:23]
  wire [31:0] mem_axi_io_axi_ar_bits_len; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_r_ready; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_r_valid; // @[SimShell.scala 39:23]
  wire [63:0] mem_axi_io_axi_r_bits_data; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_r_bits_last; // @[SimShell.scala 39:23]
  VTAMemDPI mem_dpi ( // @[SimShell.scala 38:23]
    .clock(mem_dpi_clock),
    .reset(mem_dpi_reset),
    .dpi_req_valid(mem_dpi_dpi_req_valid),
    .dpi_req_opcode(mem_dpi_dpi_req_opcode),
    .dpi_req_len(mem_dpi_dpi_req_len),
    .dpi_req_addr(mem_dpi_dpi_req_addr),
    .dpi_wr_valid(mem_dpi_dpi_wr_valid),
    .dpi_wr_bits(mem_dpi_dpi_wr_bits),
    .dpi_rd_ready(mem_dpi_dpi_rd_ready),
    .dpi_rd_valid(mem_dpi_dpi_rd_valid),
    .dpi_rd_bits(mem_dpi_dpi_rd_bits)
  );
  VTAMemDPIToAXI mem_axi ( // @[SimShell.scala 39:23]
    .clock(mem_axi_clock),
    .reset(mem_axi_reset),
    .io_dpi_req_valid(mem_axi_io_dpi_req_valid),
    .io_dpi_req_opcode(mem_axi_io_dpi_req_opcode),
    .io_dpi_req_len(mem_axi_io_dpi_req_len),
    .io_dpi_req_addr(mem_axi_io_dpi_req_addr),
    .io_dpi_wr_valid(mem_axi_io_dpi_wr_valid),
    .io_dpi_wr_bits(mem_axi_io_dpi_wr_bits),
    .io_dpi_rd_ready(mem_axi_io_dpi_rd_ready),
    .io_dpi_rd_valid(mem_axi_io_dpi_rd_valid),
    .io_dpi_rd_bits(mem_axi_io_dpi_rd_bits),
    .io_axi_aw_ready(mem_axi_io_axi_aw_ready),
    .io_axi_aw_valid(mem_axi_io_axi_aw_valid),
    .io_axi_aw_bits_addr(mem_axi_io_axi_aw_bits_addr),
    .io_axi_aw_bits_len(mem_axi_io_axi_aw_bits_len),
    .io_axi_w_ready(mem_axi_io_axi_w_ready),
    .io_axi_w_valid(mem_axi_io_axi_w_valid),
    .io_axi_w_bits_data(mem_axi_io_axi_w_bits_data),
    .io_axi_w_bits_last(mem_axi_io_axi_w_bits_last),
    .io_axi_b_ready(mem_axi_io_axi_b_ready),
    .io_axi_b_valid(mem_axi_io_axi_b_valid),
    .io_axi_ar_ready(mem_axi_io_axi_ar_ready),
    .io_axi_ar_valid(mem_axi_io_axi_ar_valid),
    .io_axi_ar_bits_addr(mem_axi_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(mem_axi_io_axi_ar_bits_len),
    .io_axi_r_ready(mem_axi_io_axi_r_ready),
    .io_axi_r_valid(mem_axi_io_axi_r_valid),
    .io_axi_r_bits_data(mem_axi_io_axi_r_bits_data),
    .io_axi_r_bits_last(mem_axi_io_axi_r_bits_last)
  );
  assign io_axi_aw_ready = mem_axi_io_axi_aw_ready; // @[SimShell.scala 43:10]
  assign io_axi_w_ready = mem_axi_io_axi_w_ready; // @[SimShell.scala 43:10]
  assign io_axi_b_valid = mem_axi_io_axi_b_valid; // @[SimShell.scala 43:10]
  assign io_axi_ar_ready = mem_axi_io_axi_ar_ready; // @[SimShell.scala 43:10]
  assign io_axi_r_valid = mem_axi_io_axi_r_valid; // @[SimShell.scala 43:10]
  assign io_axi_r_bits_data = mem_axi_io_axi_r_bits_data; // @[SimShell.scala 43:10]
  assign io_axi_r_bits_last = mem_axi_io_axi_r_bits_last; // @[SimShell.scala 43:10]
  assign mem_dpi_clock = clock; // @[SimShell.scala 41:20]
  assign mem_dpi_reset = reset; // @[SimShell.scala 40:20]
  assign mem_dpi_dpi_req_valid = mem_axi_io_dpi_req_valid; // @[SimShell.scala 42:18]
  assign mem_dpi_dpi_req_opcode = mem_axi_io_dpi_req_opcode; // @[SimShell.scala 42:18]
  assign mem_dpi_dpi_req_len = mem_axi_io_dpi_req_len; // @[SimShell.scala 42:18]
  assign mem_dpi_dpi_req_addr = mem_axi_io_dpi_req_addr; // @[SimShell.scala 42:18]
  assign mem_dpi_dpi_wr_valid = mem_axi_io_dpi_wr_valid; // @[SimShell.scala 42:18]
  assign mem_dpi_dpi_wr_bits = mem_axi_io_dpi_wr_bits; // @[SimShell.scala 42:18]
  assign mem_dpi_dpi_rd_ready = mem_axi_io_dpi_rd_ready; // @[SimShell.scala 42:18]
  assign mem_axi_clock = clock;
  assign mem_axi_reset = reset;
  assign mem_axi_io_dpi_rd_valid = mem_dpi_dpi_rd_valid; // @[SimShell.scala 42:18]
  assign mem_axi_io_dpi_rd_bits = mem_dpi_dpi_rd_bits; // @[SimShell.scala 42:18]
  assign mem_axi_io_axi_aw_valid = io_axi_aw_valid; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_aw_bits_addr = io_axi_aw_bits_addr; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_aw_bits_len = io_axi_aw_bits_len; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_w_valid = io_axi_w_valid; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_w_bits_data = io_axi_w_bits_data; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_w_bits_last = io_axi_w_bits_last; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_b_ready = io_axi_b_ready; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_ar_valid = io_axi_ar_valid; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_ar_bits_addr = io_axi_ar_bits_addr; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_ar_bits_len = io_axi_ar_bits_len; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_r_ready = io_axi_r_ready; // @[SimShell.scala 43:10]
endmodule
module AXISimShell(
  input         clock,
  input         reset,
  output        mem_aw_ready,
  input         mem_aw_valid,
  input  [31:0] mem_aw_bits_addr,
  input  [31:0] mem_aw_bits_len,
  output        mem_w_ready,
  input         mem_w_valid,
  input  [63:0] mem_w_bits_data,
  input         mem_w_bits_last,
  input         mem_b_ready,
  output        mem_b_valid,
  output        mem_ar_ready,
  input         mem_ar_valid,
  input  [31:0] mem_ar_bits_addr,
  input  [31:0] mem_ar_bits_len,
  input         mem_r_ready,
  output        mem_r_valid,
  output [63:0] mem_r_bits_data,
  output        mem_r_bits_last,
  input         host_aw_ready,
  output        host_aw_valid,
  output [31:0] host_aw_bits_addr,
  input         host_w_ready,
  output        host_w_valid,
  output [63:0] host_w_bits_data,
  output        host_b_ready,
  input         host_b_valid,
  input         host_ar_ready,
  output        host_ar_valid,
  output [31:0] host_ar_bits_addr,
  output        host_r_ready,
  input         host_r_valid,
  input  [63:0] host_r_bits_data,
  input         sim_clock,
  output        sim_wait
);
  wire  mod_sim_clock; // @[SimShell.scala 93:23]
  wire  mod_sim_reset; // @[SimShell.scala 93:23]
  wire  mod_sim_sim_wait; // @[SimShell.scala 93:23]
  wire  mod_host_clock; // @[SimShell.scala 94:24]
  wire  mod_host_reset; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_aw_ready; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_aw_valid; // @[SimShell.scala 94:24]
  wire [31:0] mod_host_io_axi_aw_bits_addr; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_w_ready; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_w_valid; // @[SimShell.scala 94:24]
  wire [63:0] mod_host_io_axi_w_bits_data; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_b_ready; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_b_valid; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_ar_ready; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_ar_valid; // @[SimShell.scala 94:24]
  wire [31:0] mod_host_io_axi_ar_bits_addr; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_r_ready; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_r_valid; // @[SimShell.scala 94:24]
  wire [63:0] mod_host_io_axi_r_bits_data; // @[SimShell.scala 94:24]
  wire  mod_mem_clock; // @[SimShell.scala 95:23]
  wire  mod_mem_reset; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_aw_ready; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_aw_valid; // @[SimShell.scala 95:23]
  wire [31:0] mod_mem_io_axi_aw_bits_addr; // @[SimShell.scala 95:23]
  wire [31:0] mod_mem_io_axi_aw_bits_len; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_w_ready; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_w_valid; // @[SimShell.scala 95:23]
  wire [63:0] mod_mem_io_axi_w_bits_data; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_w_bits_last; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_b_ready; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_b_valid; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_ar_ready; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_ar_valid; // @[SimShell.scala 95:23]
  wire [31:0] mod_mem_io_axi_ar_bits_addr; // @[SimShell.scala 95:23]
  wire [31:0] mod_mem_io_axi_ar_bits_len; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_r_ready; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_r_valid; // @[SimShell.scala 95:23]
  wire [63:0] mod_mem_io_axi_r_bits_data; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_r_bits_last; // @[SimShell.scala 95:23]
  VTASim mod_sim ( // @[SimShell.scala 93:23]
    .clock(mod_sim_clock),
    .reset(mod_sim_reset),
    .sim_wait(mod_sim_sim_wait)
  );
  VTAHost mod_host ( // @[SimShell.scala 94:24]
    .clock(mod_host_clock),
    .reset(mod_host_reset),
    .io_axi_aw_ready(mod_host_io_axi_aw_ready),
    .io_axi_aw_valid(mod_host_io_axi_aw_valid),
    .io_axi_aw_bits_addr(mod_host_io_axi_aw_bits_addr),
    .io_axi_w_ready(mod_host_io_axi_w_ready),
    .io_axi_w_valid(mod_host_io_axi_w_valid),
    .io_axi_w_bits_data(mod_host_io_axi_w_bits_data),
    .io_axi_b_ready(mod_host_io_axi_b_ready),
    .io_axi_b_valid(mod_host_io_axi_b_valid),
    .io_axi_ar_ready(mod_host_io_axi_ar_ready),
    .io_axi_ar_valid(mod_host_io_axi_ar_valid),
    .io_axi_ar_bits_addr(mod_host_io_axi_ar_bits_addr),
    .io_axi_r_ready(mod_host_io_axi_r_ready),
    .io_axi_r_valid(mod_host_io_axi_r_valid),
    .io_axi_r_bits_data(mod_host_io_axi_r_bits_data)
  );
  VTAMem mod_mem ( // @[SimShell.scala 95:23]
    .clock(mod_mem_clock),
    .reset(mod_mem_reset),
    .io_axi_aw_ready(mod_mem_io_axi_aw_ready),
    .io_axi_aw_valid(mod_mem_io_axi_aw_valid),
    .io_axi_aw_bits_addr(mod_mem_io_axi_aw_bits_addr),
    .io_axi_aw_bits_len(mod_mem_io_axi_aw_bits_len),
    .io_axi_w_ready(mod_mem_io_axi_w_ready),
    .io_axi_w_valid(mod_mem_io_axi_w_valid),
    .io_axi_w_bits_data(mod_mem_io_axi_w_bits_data),
    .io_axi_w_bits_last(mod_mem_io_axi_w_bits_last),
    .io_axi_b_ready(mod_mem_io_axi_b_ready),
    .io_axi_b_valid(mod_mem_io_axi_b_valid),
    .io_axi_ar_ready(mod_mem_io_axi_ar_ready),
    .io_axi_ar_valid(mod_mem_io_axi_ar_valid),
    .io_axi_ar_bits_addr(mod_mem_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(mod_mem_io_axi_ar_bits_len),
    .io_axi_r_ready(mod_mem_io_axi_r_ready),
    .io_axi_r_valid(mod_mem_io_axi_r_valid),
    .io_axi_r_bits_data(mod_mem_io_axi_r_bits_data),
    .io_axi_r_bits_last(mod_mem_io_axi_r_bits_last)
  );
  assign mem_aw_ready = mod_mem_io_axi_aw_ready; // @[SimShell.scala 96:7]
  assign mem_w_ready = mod_mem_io_axi_w_ready; // @[SimShell.scala 96:7]
  assign mem_b_valid = mod_mem_io_axi_b_valid; // @[SimShell.scala 96:7]
  assign mem_ar_ready = mod_mem_io_axi_ar_ready; // @[SimShell.scala 96:7]
  assign mem_r_valid = mod_mem_io_axi_r_valid; // @[SimShell.scala 96:7]
  assign mem_r_bits_data = mod_mem_io_axi_r_bits_data; // @[SimShell.scala 96:7]
  assign mem_r_bits_last = mod_mem_io_axi_r_bits_last; // @[SimShell.scala 96:7]
  assign host_aw_valid = mod_host_io_axi_aw_valid; // @[SimShell.scala 97:8]
  assign host_aw_bits_addr = mod_host_io_axi_aw_bits_addr; // @[SimShell.scala 97:8]
  assign host_w_valid = mod_host_io_axi_w_valid; // @[SimShell.scala 97:8]
  assign host_w_bits_data = mod_host_io_axi_w_bits_data; // @[SimShell.scala 97:8]
  assign host_b_ready = mod_host_io_axi_b_ready; // @[SimShell.scala 97:8]
  assign host_ar_valid = mod_host_io_axi_ar_valid; // @[SimShell.scala 97:8]
  assign host_ar_bits_addr = mod_host_io_axi_ar_bits_addr; // @[SimShell.scala 97:8]
  assign host_r_ready = mod_host_io_axi_r_ready; // @[SimShell.scala 97:8]
  assign sim_wait = mod_sim_sim_wait; // @[SimShell.scala 100:12]
  assign mod_sim_clock = sim_clock; // @[SimShell.scala 99:17]
  assign mod_sim_reset = reset; // @[SimShell.scala 98:17]
  assign mod_host_clock = clock;
  assign mod_host_reset = reset;
  assign mod_host_io_axi_aw_ready = host_aw_ready; // @[SimShell.scala 97:8]
  assign mod_host_io_axi_w_ready = host_w_ready; // @[SimShell.scala 97:8]
  assign mod_host_io_axi_b_valid = host_b_valid; // @[SimShell.scala 97:8]
  assign mod_host_io_axi_ar_ready = host_ar_ready; // @[SimShell.scala 97:8]
  assign mod_host_io_axi_r_valid = host_r_valid; // @[SimShell.scala 97:8]
  assign mod_host_io_axi_r_bits_data = host_r_bits_data; // @[SimShell.scala 97:8]
  assign mod_mem_clock = clock;
  assign mod_mem_reset = reset;
  assign mod_mem_io_axi_aw_valid = mem_aw_valid; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_aw_bits_addr = mem_aw_bits_addr; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_aw_bits_len = mem_aw_bits_len; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_w_valid = mem_w_valid; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_w_bits_data = mem_w_bits_data; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_w_bits_last = mem_w_bits_last; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_b_ready = mem_b_ready; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_ar_valid = mem_ar_valid; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_ar_bits_addr = mem_ar_bits_addr; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_ar_bits_len = mem_ar_bits_len; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_r_ready = mem_r_ready; // @[SimShell.scala 96:7]
endmodule
module DCR(
  input         clock,
  input         reset,
  output        io_host_aw_ready,
  input         io_host_aw_valid,
  input  [31:0] io_host_aw_bits_addr,
  output        io_host_w_ready,
  input         io_host_w_valid,
  input  [63:0] io_host_w_bits_data,
  input         io_host_b_ready,
  output        io_host_b_valid,
  output        io_host_ar_ready,
  input         io_host_ar_valid,
  input  [31:0] io_host_ar_bits_addr,
  input         io_host_r_ready,
  output        io_host_r_valid,
  output [63:0] io_host_r_bits_data,
  output        io_dcr_launch,
  input         io_dcr_finish,
  input         io_dcr_ecnt_0_valid,
  input  [31:0] io_dcr_ecnt_0_bits,
  input  [31:0] io_dcr_ecnt_1_bits,
  input  [31:0] io_dcr_ecnt_2_bits,
  input  [31:0] io_dcr_ecnt_3_bits,
  input  [31:0] io_dcr_ecnt_4_bits,
  input  [31:0] io_dcr_ecnt_5_bits,
  input  [31:0] io_dcr_ecnt_6_bits,
  output [31:0] io_dcr_vals_0,
  output [31:0] io_dcr_ptrs_0,
  output [31:0] io_dcr_ptrs_1,
  output [31:0] io_dcr_ptrs_2,
  output [31:0] io_dcr_ptrs_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] waddr; // @[DCR.scala 88:22]
  reg [1:0] wstate; // @[DCR.scala 91:23]
  reg  rstate; // @[DCR.scala 95:23]
  reg [31:0] rdata; // @[DCR.scala 96:22]
  reg [31:0] reg_0; // @[DCR.scala 102:37]
  reg [31:0] reg_1; // @[DCR.scala 102:37]
  reg [31:0] reg_2; // @[DCR.scala 102:37]
  reg [31:0] reg_3; // @[DCR.scala 102:37]
  reg [31:0] reg_4; // @[DCR.scala 102:37]
  reg [31:0] reg_5; // @[DCR.scala 102:37]
  reg [31:0] reg_6; // @[DCR.scala 102:37]
  reg [31:0] reg_7; // @[DCR.scala 102:37]
  reg [31:0] reg_18; // @[DCR.scala 102:37]
  reg [31:0] reg_19; // @[DCR.scala 102:37]
  reg [31:0] reg_20; // @[DCR.scala 102:37]
  reg [31:0] reg_21; // @[DCR.scala 102:37]
  reg [31:0] reg_22; // @[DCR.scala 102:37]
  wire  _T = 2'h0 == wstate; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == wstate; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h2 == wstate; // @[Conditional.scala 37:30]
  wire  _T_3 = io_host_aw_ready & io_host_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_7 = ~rstate; // @[Conditional.scala 37:30]
  wire  _GEN_7 = io_host_ar_valid | rstate; // @[DCR.scala 138:30]
  wire  _T_11 = io_host_w_ready & io_host_w_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = 32'h0 == waddr; // @[DCR.scala 156:44]
  wire  _T_13 = _T_11 & _T_12; // @[DCR.scala 156:31]
  wire [63:0] _GEN_11 = _T_13 ? io_host_w_bits_data : {{32'd0}, reg_0}; // @[DCR.scala 156:55]
  wire [63:0] _GEN_12 = io_dcr_finish ? 64'h2 : _GEN_11; // @[DCR.scala 154:23]
  wire  _T_15 = 32'h4 == waddr; // @[DCR.scala 163:51]
  wire  _T_16 = _T_11 & _T_15; // @[DCR.scala 163:33]
  wire [63:0] _GEN_13 = _T_16 ? io_host_w_bits_data : {{32'd0}, reg_1}; // @[DCR.scala 163:62]
  wire [63:0] _GEN_14 = io_dcr_ecnt_0_valid ? {{32'd0}, io_dcr_ecnt_0_bits} : _GEN_13; // @[DCR.scala 161:32]
  wire [63:0] _GEN_16 = {{32'd0}, io_dcr_ecnt_1_bits}; // @[DCR.scala 161:32]
  wire [63:0] _GEN_18 = {{32'd0}, io_dcr_ecnt_2_bits}; // @[DCR.scala 161:32]
  wire [63:0] _GEN_20 = {{32'd0}, io_dcr_ecnt_3_bits}; // @[DCR.scala 161:32]
  wire [63:0] _GEN_22 = {{32'd0}, io_dcr_ecnt_4_bits}; // @[DCR.scala 161:32]
  wire [63:0] _GEN_24 = {{32'd0}, io_dcr_ecnt_5_bits}; // @[DCR.scala 161:32]
  wire [63:0] _GEN_26 = {{32'd0}, io_dcr_ecnt_6_bits}; // @[DCR.scala 161:32]
  wire  _T_66 = 32'h48 == waddr; // @[DCR.scala 169:45]
  wire  _T_67 = _T_11 & _T_66; // @[DCR.scala 169:27]
  wire [63:0] _GEN_47 = _T_67 ? io_host_w_bits_data : {{32'd0}, reg_18}; // @[DCR.scala 169:56]
  wire  _T_69 = 32'h4c == waddr; // @[DCR.scala 169:45]
  wire  _T_70 = _T_11 & _T_69; // @[DCR.scala 169:27]
  wire [63:0] _GEN_48 = _T_70 ? io_host_w_bits_data : {{32'd0}, reg_19}; // @[DCR.scala 169:56]
  wire  _T_72 = 32'h50 == waddr; // @[DCR.scala 169:45]
  wire  _T_73 = _T_11 & _T_72; // @[DCR.scala 169:27]
  wire [63:0] _GEN_49 = _T_73 ? io_host_w_bits_data : {{32'd0}, reg_20}; // @[DCR.scala 169:56]
  wire  _T_75 = 32'h54 == waddr; // @[DCR.scala 169:45]
  wire  _T_76 = _T_11 & _T_75; // @[DCR.scala 169:27]
  wire [63:0] _GEN_50 = _T_76 ? io_host_w_bits_data : {{32'd0}, reg_21}; // @[DCR.scala 169:56]
  wire  _T_78 = 32'h58 == waddr; // @[DCR.scala 169:45]
  wire  _T_79 = _T_11 & _T_78; // @[DCR.scala 169:27]
  wire [63:0] _GEN_51 = _T_79 ? io_host_w_bits_data : {{32'd0}, reg_22}; // @[DCR.scala 169:56]
  wire  _T_80 = io_host_ar_ready & io_host_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_81 = 32'h0 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_83 = 32'h4 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_85 = 32'h8 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_87 = 32'hc == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_89 = 32'h10 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_91 = 32'h14 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_93 = 32'h18 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_95 = 32'h1c == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_97 = 32'h20 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_99 = 32'h24 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_101 = 32'h28 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_103 = 32'h2c == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_105 = 32'h30 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_107 = 32'h34 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_109 = 32'h38 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_111 = 32'h3c == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_113 = 32'h40 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_115 = 32'h44 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_117 = 32'h48 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_119 = 32'h4c == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_121 = 32'h50 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_123 = 32'h54 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_125 = 32'h58 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  assign io_host_aw_ready = wstate == 2'h0; // @[DCR.scala 131:20]
  assign io_host_w_ready = wstate == 2'h1; // @[DCR.scala 132:19]
  assign io_host_b_valid = wstate == 2'h2; // @[DCR.scala 133:19]
  assign io_host_ar_ready = ~rstate; // @[DCR.scala 149:20]
  assign io_host_r_valid = rstate; // @[DCR.scala 150:19]
  assign io_host_r_bits_data = {{32'd0}, rdata}; // @[DCR.scala 151:23]
  assign io_dcr_launch = reg_0[0]; // @[DCR.scala 178:17]
  assign io_dcr_vals_0 = reg_18; // @[DCR.scala 181:20]
  assign io_dcr_ptrs_0 = reg_19; // @[DCR.scala 186:22]
  assign io_dcr_ptrs_1 = reg_20; // @[DCR.scala 186:22]
  assign io_dcr_ptrs_2 = reg_21; // @[DCR.scala 186:22]
  assign io_dcr_ptrs_3 = reg_22; // @[DCR.scala 186:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waddr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  wstate = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  rstate = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  rdata = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_0 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_4 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_5 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_6 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_7 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_18 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_19 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_20 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_21 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_22 = _RAND_16[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      waddr <= 32'hffff;
    end else if (_T_3) begin
      waddr <= io_host_aw_bits_addr;
    end
    if (reset) begin
      wstate <= 2'h0;
    end else if (_T) begin
      if (io_host_aw_valid) begin
        wstate <= 2'h1;
      end
    end else if (_T_1) begin
      if (io_host_w_valid) begin
        wstate <= 2'h2;
      end
    end else if (_T_2) begin
      if (io_host_b_ready) begin
        wstate <= 2'h0;
      end
    end
    if (reset) begin
      rstate <= 1'h0;
    end else if (_T_7) begin
      rstate <= _GEN_7;
    end else if (rstate) begin
      if (io_host_r_ready) begin
        rstate <= 1'h0;
      end
    end
    if (reset) begin
      rdata <= 32'h0;
    end else if (_T_80) begin
      if (_T_125) begin
        rdata <= reg_22;
      end else if (_T_123) begin
        rdata <= reg_21;
      end else if (_T_121) begin
        rdata <= reg_20;
      end else if (_T_119) begin
        rdata <= reg_19;
      end else if (_T_117) begin
        rdata <= reg_18;
      end else if (_T_115) begin
        rdata <= 32'h0;
      end else if (_T_113) begin
        rdata <= 32'h0;
      end else if (_T_111) begin
        rdata <= 32'h0;
      end else if (_T_109) begin
        rdata <= 32'h0;
      end else if (_T_107) begin
        rdata <= 32'h0;
      end else if (_T_105) begin
        rdata <= 32'h0;
      end else if (_T_103) begin
        rdata <= 32'h0;
      end else if (_T_101) begin
        rdata <= 32'h0;
      end else if (_T_99) begin
        rdata <= 32'h0;
      end else if (_T_97) begin
        rdata <= 32'h0;
      end else if (_T_95) begin
        rdata <= reg_7;
      end else if (_T_93) begin
        rdata <= reg_6;
      end else if (_T_91) begin
        rdata <= reg_5;
      end else if (_T_89) begin
        rdata <= reg_4;
      end else if (_T_87) begin
        rdata <= reg_3;
      end else if (_T_85) begin
        rdata <= reg_2;
      end else if (_T_83) begin
        rdata <= reg_1;
      end else if (_T_81) begin
        rdata <= reg_0;
      end else begin
        rdata <= 32'h0;
      end
    end
    if (reset) begin
      reg_0 <= 32'h0;
    end else begin
      reg_0 <= _GEN_12[31:0];
    end
    if (reset) begin
      reg_1 <= 32'h0;
    end else begin
      reg_1 <= _GEN_14[31:0];
    end
    if (reset) begin
      reg_2 <= 32'h0;
    end else begin
      reg_2 <= _GEN_16[31:0];
    end
    if (reset) begin
      reg_3 <= 32'h0;
    end else begin
      reg_3 <= _GEN_18[31:0];
    end
    if (reset) begin
      reg_4 <= 32'h0;
    end else begin
      reg_4 <= _GEN_20[31:0];
    end
    if (reset) begin
      reg_5 <= 32'h0;
    end else begin
      reg_5 <= _GEN_22[31:0];
    end
    if (reset) begin
      reg_6 <= 32'h0;
    end else begin
      reg_6 <= _GEN_24[31:0];
    end
    if (reset) begin
      reg_7 <= 32'h0;
    end else begin
      reg_7 <= _GEN_26[31:0];
    end
    if (reset) begin
      reg_18 <= 32'h0;
    end else begin
      reg_18 <= _GEN_47[31:0];
    end
    if (reset) begin
      reg_19 <= 32'h0;
    end else begin
      reg_19 <= _GEN_48[31:0];
    end
    if (reset) begin
      reg_20 <= 32'h0;
    end else begin
      reg_20 <= _GEN_49[31:0];
    end
    if (reset) begin
      reg_21 <= 32'h0;
    end else begin
      reg_21 <= _GEN_50[31:0];
    end
    if (reset) begin
      reg_22 <= 32'h0;
    end else begin
      reg_22 <= _GEN_51[31:0];
    end
  end
endmodule
module Arbiter(
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [1:0]  io_chosen
);
  wire [1:0] _GEN_0 = io_in_1_valid ? 2'h1 : 2'h2; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_2 = io_in_1_valid ? io_in_1_bits_addr : io_in_2_bits_addr; // @[Arbiter.scala 126:27]
  wire  _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  grant_2 = ~_T; // @[Arbiter.scala 31:78]
  wire  _T_4 = ~grant_2; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_4 | io_in_2_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_2; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_chosen = io_in_0_valid ? 2'h0 : _GEN_0; // @[Arbiter.scala 123:13 Arbiter.scala 127:17 Arbiter.scala 127:17]
endmodule
module DME(
  input         clock,
  input         reset,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output        io_mem_w_bits_last,
  output        io_mem_b_ready,
  input         io_mem_b_valid,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last,
  input         io_dme_rd_0_cmd_valid,
  input  [31:0] io_dme_rd_0_cmd_bits_addr,
  input         io_dme_rd_0_data_ready,
  output        io_dme_rd_0_data_valid,
  output [63:0] io_dme_rd_0_data_bits,
  input         io_dme_rd_1_cmd_valid,
  input  [31:0] io_dme_rd_1_cmd_bits_addr,
  input         io_dme_rd_1_data_ready,
  output        io_dme_rd_1_data_valid,
  output [63:0] io_dme_rd_1_data_bits,
  input         io_dme_rd_2_cmd_valid,
  input  [31:0] io_dme_rd_2_cmd_bits_addr,
  input         io_dme_rd_2_data_ready,
  output        io_dme_rd_2_data_valid,
  output [63:0] io_dme_rd_2_data_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  rd_arb_io_in_0_valid; // @[DME.scala 130:22]
  wire [31:0] rd_arb_io_in_0_bits_addr; // @[DME.scala 130:22]
  wire  rd_arb_io_in_1_valid; // @[DME.scala 130:22]
  wire [31:0] rd_arb_io_in_1_bits_addr; // @[DME.scala 130:22]
  wire  rd_arb_io_in_2_valid; // @[DME.scala 130:22]
  wire [31:0] rd_arb_io_in_2_bits_addr; // @[DME.scala 130:22]
  wire  rd_arb_io_out_ready; // @[DME.scala 130:22]
  wire  rd_arb_io_out_valid; // @[DME.scala 130:22]
  wire [31:0] rd_arb_io_out_bits_addr; // @[DME.scala 130:22]
  wire [1:0] rd_arb_io_chosen; // @[DME.scala 130:22]
  wire  _T = rd_arb_io_out_ready & rd_arb_io_out_valid; // @[Decoupled.scala 40:37]
  reg [1:0] rd_arb_chosen; // @[Reg.scala 15:16]
  reg [1:0] rstate; // @[DME.scala 138:23]
  wire  _T_1 = 2'h0 == rstate; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h1 == rstate; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h2 == rstate; // @[Conditional.scala 37:30]
  wire  _T_4 = io_mem_r_ready & io_mem_r_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = _T_4 & io_mem_r_bits_last; // @[DME.scala 152:28]
  reg [1:0] wstate; // @[DME.scala 168:23]
  reg [31:0] wr_cnt; // @[DME.scala 171:23]
  wire  _T_7 = wstate == 2'h0; // @[DME.scala 174:15]
  wire  _T_8 = io_mem_w_ready & io_mem_w_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _T_10 = wr_cnt + 32'h1; // @[DME.scala 177:22]
  wire  _T_11 = 2'h0 == wstate; // @[Conditional.scala 37:30]
  wire  _T_12 = 2'h1 == wstate; // @[Conditional.scala 37:30]
  wire  _T_13 = 2'h2 == wstate; // @[Conditional.scala 37:30]
  wire  _T_17 = 2'h3 == wstate; // @[Conditional.scala 37:30]
  reg [31:0] rd_addr; // @[Reg.scala 27:20]
  wire  _T_24 = rd_arb_chosen == 2'h0; // @[DME.scala 215:46]
  wire  _T_26 = rd_arb_chosen == 2'h1; // @[DME.scala 215:46]
  wire  _T_28 = rd_arb_chosen == 2'h2; // @[DME.scala 215:46]
  wire  _T_43 = rstate == 2'h2; // @[DME.scala 240:28]
  wire  _GEN_33 = 2'h1 == rd_arb_chosen ? io_dme_rd_1_data_ready : io_dme_rd_0_data_ready; // @[DME.scala 240:42]
  wire  _GEN_40 = 2'h2 == rd_arb_chosen ? io_dme_rd_2_data_ready : _GEN_33; // @[DME.scala 240:42]
  Arbiter rd_arb ( // @[DME.scala 130:22]
    .io_in_0_valid(rd_arb_io_in_0_valid),
    .io_in_0_bits_addr(rd_arb_io_in_0_bits_addr),
    .io_in_1_valid(rd_arb_io_in_1_valid),
    .io_in_1_bits_addr(rd_arb_io_in_1_bits_addr),
    .io_in_2_valid(rd_arb_io_in_2_valid),
    .io_in_2_bits_addr(rd_arb_io_in_2_bits_addr),
    .io_out_ready(rd_arb_io_out_ready),
    .io_out_valid(rd_arb_io_out_valid),
    .io_out_bits_addr(rd_arb_io_out_bits_addr),
    .io_chosen(rd_arb_io_chosen)
  );
  assign io_mem_aw_valid = wstate == 2'h1; // @[DME.scala 226:19]
  assign io_mem_w_valid = 1'h0; // @[DME.scala 230:18]
  assign io_mem_w_bits_last = wr_cnt == 32'h0; // @[DME.scala 232:22]
  assign io_mem_b_ready = wstate == 2'h3; // @[DME.scala 234:18]
  assign io_mem_ar_valid = rstate == 2'h1; // @[DME.scala 236:19]
  assign io_mem_ar_bits_addr = rd_addr; // @[DME.scala 237:23]
  assign io_mem_r_ready = _T_43 & _GEN_40; // @[DME.scala 240:18]
  assign io_dme_rd_0_data_valid = _T_24 & io_mem_r_valid; // @[DME.scala 215:29]
  assign io_dme_rd_0_data_bits = io_mem_r_bits_data; // @[DME.scala 216:28]
  assign io_dme_rd_1_data_valid = _T_26 & io_mem_r_valid; // @[DME.scala 215:29]
  assign io_dme_rd_1_data_bits = io_mem_r_bits_data; // @[DME.scala 216:28]
  assign io_dme_rd_2_data_valid = _T_28 & io_mem_r_valid; // @[DME.scala 215:29]
  assign io_dme_rd_2_data_bits = io_mem_r_bits_data; // @[DME.scala 216:28]
  assign rd_arb_io_in_0_valid = io_dme_rd_0_cmd_valid; // @[DME.scala 134:21]
  assign rd_arb_io_in_0_bits_addr = io_dme_rd_0_cmd_bits_addr; // @[DME.scala 134:21]
  assign rd_arb_io_in_1_valid = io_dme_rd_1_cmd_valid; // @[DME.scala 134:21]
  assign rd_arb_io_in_1_bits_addr = io_dme_rd_1_cmd_bits_addr; // @[DME.scala 134:21]
  assign rd_arb_io_in_2_valid = io_dme_rd_2_cmd_valid; // @[DME.scala 134:21]
  assign rd_arb_io_in_2_bits_addr = io_dme_rd_2_cmd_bits_addr; // @[DME.scala 134:21]
  assign rd_arb_io_out_ready = rstate == 2'h0; // @[DME.scala 210:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rd_arb_chosen = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  rstate = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  wstate = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  wr_cnt = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  rd_addr = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T) begin
      rd_arb_chosen <= rd_arb_io_chosen;
    end
    if (reset) begin
      rstate <= 2'h0;
    end else if (_T_1) begin
      if (rd_arb_io_out_valid) begin
        rstate <= 2'h1;
      end
    end else if (_T_2) begin
      if (io_mem_ar_ready) begin
        rstate <= 2'h2;
      end
    end else if (_T_3) begin
      if (_T_5) begin
        rstate <= 2'h0;
      end
    end
    if (reset) begin
      wstate <= 2'h0;
    end else if (!(_T_11)) begin
      if (_T_12) begin
        if (io_mem_aw_ready) begin
          wstate <= 2'h2;
        end
      end else if (!(_T_13)) begin
        if (_T_17) begin
          if (io_mem_b_valid) begin
            wstate <= 2'h0;
          end
        end
      end
    end
    if (reset) begin
      wr_cnt <= 32'h0;
    end else if (_T_7) begin
      wr_cnt <= 32'h0;
    end else if (_T_8) begin
      wr_cnt <= _T_10;
    end
    if (reset) begin
      rd_addr <= 32'h0;
    end else if (_T) begin
      rd_addr <= rd_arb_io_out_bits_addr;
    end
  end
endmodule
module memoryWrapper(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [7:0]  io_in_bits_inst,
  input  [63:0] io_in_bits_data,
  input  [2:0]  io_in_bits_src,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output        io_mem_b_ready,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [15:0] io_mem_ar_bits_len,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [63:0] io_out_bits_data,
  output [2:0]  io_out_bits_dst
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] addrReg; // @[mainMemWrapper.scala 36:26]
  reg [2:0] numberOfLines; // @[mainMemWrapper.scala 37:32]
  reg [2:0] srcReg; // @[mainMemWrapper.scala 38:25]
  reg [31:0] returnAddr; // @[mainMemWrapper.scala 39:29]
  reg [63:0] dataRegRead_0; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegRead_1; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegRead_2; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegRead_3; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegRead_4; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegRead_5; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegRead_6; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegWrite_0; // @[mainMemWrapper.scala 41:31]
  reg [2:0] stReg; // @[mainMemWrapper.scala 44:24]
  wire  _T_2 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = stReg == 3'h0; // @[mainMemWrapper.scala 47:35]
  wire  _T_4 = _T_2 & _T_3; // @[mainMemWrapper.scala 47:27]
  wire  _T_6 = io_in_bits_data[31:0] != 32'h0; // @[mainMemWrapper.scala 47:80]
  wire  start = _T_4 & _T_6; // @[mainMemWrapper.scala 47:46]
  wire [31:0] _T_9 = {io_in_bits_data[31:3], 3'h0}; // @[mainMemWrapper.scala 50:58]
  wire  _T_11 = io_in_bits_data[2:0] == 3'h0; // @[mainMemWrapper.scala 51:51]
  wire  _T_15 = io_in_bits_inst == 8'h1; // @[mainMemWrapper.scala 58:54]
  wire  writeInst = start & _T_15; // @[mainMemWrapper.scala 58:36]
  wire  _T_17 = io_mem_r_ready & io_mem_r_valid; // @[Decoupled.scala 40:37]
  reg [2:0] readCount; // @[Counter.scala 29:33]
  wire  _T_18 = readCount == 3'h6; // @[Counter.scala 38:24]
  wire [2:0] _T_20 = readCount + 3'h1; // @[Counter.scala 39:22]
  wire  writeWrapped = io_mem_w_ready & io_mem_w_valid; // @[Decoupled.scala 40:37]
  wire  _T_22 = stReg == 3'h5; // @[mainMemWrapper.scala 65:55]
  reg [19:0] dramLatencyCnt; // @[Counter.scala 29:33]
  wire  _T_24 = dramLatencyCnt == 20'hf423f; // @[Counter.scala 38:24]
  wire [19:0] _T_26 = dramLatencyCnt + 20'h1; // @[Counter.scala 39:22]
  wire  _T_27 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [19:0] nextPacket; // @[Counter.scala 29:33]
  wire  _T_29 = nextPacket == 20'hf423f; // @[Counter.scala 38:24]
  wire [19:0] _T_31 = nextPacket + 20'h1; // @[Counter.scala 39:22]
  wire [2:0] _T_33 = numberOfLines - 3'h1; // @[mainMemWrapper.scala 67:62]
  wire [19:0] _GEN_75 = {{17'd0}, _T_33}; // @[mainMemWrapper.scala 67:44]
  wire  packetsDone = nextPacket == _GEN_75; // @[mainMemWrapper.scala 67:44]
  wire [31:0] _T_38 = returnAddr + 32'h8; // @[mainMemWrapper.scala 70:34]
  wire  _T_43 = stReg == 3'h1; // @[mainMemWrapper.scala 82:38]
  wire  _T_45 = stReg == 3'h2; // @[mainMemWrapper.scala 85:37]
  wire [3:0] _T_47 = 3'h1 * numberOfLines; // @[mainMemWrapper.scala 89:35]
  wire [3:0] _T_49 = _T_47 - 4'h1; // @[mainMemWrapper.scala 89:51]
  wire [20:0] _T_51 = nextPacket * 20'h1; // @[mainMemWrapper.scala 101:78]
  wire [21:0] _T_52 = {{1'd0}, _T_51}; // @[mainMemWrapper.scala 101:88]
  wire [63:0] _GEN_34 = 3'h1 == _T_52[2:0] ? dataRegRead_1 : dataRegRead_0; // @[mainMemWrapper.scala 101:22]
  wire [63:0] _GEN_35 = 3'h2 == _T_52[2:0] ? dataRegRead_2 : _GEN_34; // @[mainMemWrapper.scala 101:22]
  wire [63:0] _GEN_36 = 3'h3 == _T_52[2:0] ? dataRegRead_3 : _GEN_35; // @[mainMemWrapper.scala 101:22]
  wire [63:0] _GEN_37 = 3'h4 == _T_52[2:0] ? dataRegRead_4 : _GEN_36; // @[mainMemWrapper.scala 101:22]
  wire [63:0] _GEN_38 = 3'h5 == _T_52[2:0] ? dataRegRead_5 : _GEN_37; // @[mainMemWrapper.scala 101:22]
  wire  _T_55 = 3'h0 == stReg; // @[Conditional.scala 37:30]
  wire  _T_56 = 3'h3 == stReg; // @[Conditional.scala 37:30]
  wire  _T_57 = io_mem_ar_ready & io_mem_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_58 = 3'h4 == stReg; // @[Conditional.scala 37:30]
  wire  _T_60 = _T_17 & io_mem_r_bits_last; // @[mainMemWrapper.scala 129:34]
  wire  _T_61 = 3'h1 == stReg; // @[Conditional.scala 37:30]
  wire  _T_62 = io_mem_aw_ready & io_mem_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_63 = 3'h2 == stReg; // @[Conditional.scala 37:30]
  wire  _T_64 = 3'h5 == stReg; // @[Conditional.scala 37:30]
  wire  _T_65 = dramLatencyCnt > 20'hc8; // @[mainMemWrapper.scala 146:34]
  wire  _T_67 = packetsDone & _T_27; // @[mainMemWrapper.scala 148:34]
  wire  _GEN_49 = _T_64 & _T_65; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_63 ? 1'h0 : _GEN_49; // @[Conditional.scala 39:67]
  wire  _GEN_56 = _T_61 ? 1'h0 : _T_63; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_61 ? 1'h0 : _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_60 = _T_58 ? 1'h0 : _T_61; // @[Conditional.scala 39:67]
  wire  _GEN_61 = _T_58 ? 1'h0 : _GEN_56; // @[Conditional.scala 39:67]
  wire  _GEN_62 = _T_58 ? 1'h0 : _GEN_57; // @[Conditional.scala 39:67]
  wire  _GEN_65 = _T_56 ? 1'h0 : _T_58; // @[Conditional.scala 39:67]
  wire  _GEN_66 = _T_56 ? 1'h0 : _GEN_60; // @[Conditional.scala 39:67]
  wire  _GEN_67 = _T_56 ? 1'h0 : _GEN_61; // @[Conditional.scala 39:67]
  wire  _GEN_68 = _T_56 ? 1'h0 : _GEN_62; // @[Conditional.scala 39:67]
  assign io_in_ready = stReg == 3'h0; // @[mainMemWrapper.scala 56:17]
  assign io_mem_aw_valid = _T_55 ? 1'h0 : _GEN_66; // @[mainMemWrapper.scala 93:21 mainMemWrapper.scala 134:29]
  assign io_mem_aw_bits_addr = _T_43 ? addrReg : 32'h0; // @[mainMemWrapper.scala 82:25]
  assign io_mem_w_valid = _T_55 ? 1'h0 : _GEN_67; // @[mainMemWrapper.scala 95:20 mainMemWrapper.scala 140:28]
  assign io_mem_w_bits_data = _T_45 ? dataRegWrite_0 : 64'h0; // @[mainMemWrapper.scala 85:24]
  assign io_mem_b_ready = stReg == 3'h2; // @[mainMemWrapper.scala 90:20]
  assign io_mem_ar_valid = _T_55 ? 1'h0 : _T_56; // @[mainMemWrapper.scala 92:21 mainMemWrapper.scala 122:29]
  assign io_mem_ar_bits_addr = addrReg; // @[mainMemWrapper.scala 88:25]
  assign io_mem_ar_bits_len = {{12'd0}, _T_49}; // @[mainMemWrapper.scala 89:24]
  assign io_mem_r_ready = _T_55 ? 1'h0 : _GEN_65; // @[mainMemWrapper.scala 94:20 mainMemWrapper.scala 128:28]
  assign io_out_valid = _T_55 ? 1'h0 : _GEN_68; // @[mainMemWrapper.scala 109:18 mainMemWrapper.scala 147:30]
  assign io_out_bits_addr = returnAddr; // @[mainMemWrapper.scala 102:22]
  assign io_out_bits_data = 3'h6 == _T_52[2:0] ? dataRegRead_6 : _GEN_38; // @[mainMemWrapper.scala 101:22]
  assign io_out_bits_dst = srcReg; // @[mainMemWrapper.scala 105:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addrReg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  numberOfLines = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  srcReg = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  returnAddr = _RAND_3[31:0];
  _RAND_4 = {2{`RANDOM}};
  dataRegRead_0 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  dataRegRead_1 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataRegRead_2 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataRegRead_3 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataRegRead_4 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  dataRegRead_5 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  dataRegRead_6 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  dataRegWrite_0 = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  stReg = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  readCount = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  dramLatencyCnt = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  nextPacket = _RAND_15[19:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addrReg <= 32'h0;
    end else if (start) begin
      addrReg <= _T_9;
    end
    if (reset) begin
      numberOfLines <= 3'h0;
    end else if (start) begin
      if (_T_11) begin
        numberOfLines <= 3'h1;
      end else begin
        numberOfLines <= io_in_bits_data[2:0];
      end
    end
    if (reset) begin
      srcReg <= 3'h0;
    end else if (start) begin
      srcReg <= io_in_bits_src;
    end
    if (reset) begin
      returnAddr <= 32'h0;
    end else if (_T_27) begin
      returnAddr <= _T_38;
    end else if (start) begin
      returnAddr <= io_in_bits_addr;
    end
    if (reset) begin
      dataRegRead_0 <= 64'h0;
    end else if (_T_17) begin
      if (3'h0 == readCount) begin
        dataRegRead_0 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegRead_1 <= 64'h0;
    end else if (_T_17) begin
      if (3'h1 == readCount) begin
        dataRegRead_1 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegRead_2 <= 64'h0;
    end else if (_T_17) begin
      if (3'h2 == readCount) begin
        dataRegRead_2 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegRead_3 <= 64'h0;
    end else if (_T_17) begin
      if (3'h3 == readCount) begin
        dataRegRead_3 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegRead_4 <= 64'h0;
    end else if (_T_17) begin
      if (3'h4 == readCount) begin
        dataRegRead_4 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegRead_5 <= 64'h0;
    end else if (_T_17) begin
      if (3'h5 == readCount) begin
        dataRegRead_5 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegRead_6 <= 64'h0;
    end else if (_T_17) begin
      if (3'h6 == readCount) begin
        dataRegRead_6 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegWrite_0 <= 64'h0;
    end else if (writeInst) begin
      dataRegWrite_0 <= io_in_bits_data;
    end
    if (reset) begin
      stReg <= 3'h0;
    end else if (_T_55) begin
      if (start) begin
        if (writeInst) begin
          stReg <= 3'h1;
        end else begin
          stReg <= 3'h3;
        end
      end
    end else if (_T_56) begin
      if (_T_57) begin
        stReg <= 3'h4;
      end
    end else if (_T_58) begin
      if (_T_60) begin
        stReg <= 3'h5;
      end
    end else if (_T_61) begin
      if (_T_62) begin
        stReg <= 3'h2;
      end
    end else if (_T_63) begin
      if (writeWrapped) begin
        stReg <= 3'h0;
      end
    end else if (_T_64) begin
      if (_T_65) begin
        if (_T_67) begin
          stReg <= 3'h0;
        end
      end
    end
    if (reset) begin
      readCount <= 3'h0;
    end else if (start) begin
      readCount <= 3'h0;
    end else if (_T_17) begin
      if (_T_18) begin
        readCount <= 3'h0;
      end else begin
        readCount <= _T_20;
      end
    end
    if (reset) begin
      dramLatencyCnt <= 20'h0;
    end else if (start) begin
      dramLatencyCnt <= 20'h0;
    end else if (_T_22) begin
      if (_T_24) begin
        dramLatencyCnt <= 20'h0;
      end else begin
        dramLatencyCnt <= _T_26;
      end
    end
    if (reset) begin
      nextPacket <= 20'h0;
    end else if (start) begin
      nextPacket <= 20'h0;
    end else if (_T_27) begin
      if (_T_29) begin
        nextPacket <= 20'h0;
      end else begin
        nextPacket <= _T_31;
      end
    end
  end
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_inst,
  input  [63:0] io_enq_bits_data,
  input  [2:0]  io_enq_bits_src,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_inst,
  output [63:0] io_deq_bits_data,
  output [2:0]  io_deq_bits_src
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:0]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_7_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [7:0] ram_inst [0:0]; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_7_addr; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:0]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_7_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_src [0:0]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_src__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_src__T_7_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_src__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_en; // @[Decoupled.scala 209:16]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram_addr__T_7_addr = 1'h0;
  assign ram_addr__T_7_data = ram_addr[ram_addr__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_3_data = io_enq_bits_addr;
  assign ram_addr__T_3_addr = 1'h0;
  assign ram_addr__T_3_mask = 1'h1;
  assign ram_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst__T_7_addr = 1'h0;
  assign ram_inst__T_7_data = ram_inst[ram_inst__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst__T_3_data = io_enq_bits_inst;
  assign ram_inst__T_3_addr = 1'h0;
  assign ram_inst__T_3_mask = 1'h1;
  assign ram_inst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_7_addr = 1'h0;
  assign ram_data__T_7_data = ram_data[ram_data__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = 1'h0;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_src__T_7_addr = 1'h0;
  assign ram_src__T_7_data = ram_src[ram_src__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_src__T_3_data = io_enq_bits_src;
  assign ram_src__T_3_addr = 1'h0;
  assign ram_src__T_3_mask = 1'h1;
  assign ram_src__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst = ram_inst__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_src = ram_src__T_7_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_inst[initvar] = _RAND_1[7:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_src[initvar] = _RAND_3[2:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_3_en & ram_addr__T_3_mask) begin
      ram_addr[ram_addr__T_3_addr] <= ram_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst__T_3_en & ram_inst__T_3_mask) begin
      ram_inst[ram_inst__T_3_addr] <= ram_inst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_src__T_3_en & ram_src__T_3_mask) begin
      ram_src[ram_src__T_3_addr] <= ram_src__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_4) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_inst,
  input  [63:0] io_enq_bits_data,
  input  [2:0]  io_enq_bits_src,
  input  [2:0]  io_enq_bits_dst,
  input  [1:0]  io_enq_bits_msgType,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_inst,
  output [63:0] io_deq_bits_data,
  output [2:0]  io_deq_bits_src,
  output [2:0]  io_deq_bits_dst,
  output [1:0]  io_deq_bits_msgType
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:1]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_11_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [7:0] ram_inst [0:1]; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_11_addr; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_11_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_src [0:1]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_src__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_src__T_11_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_src__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_dst [0:1]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_dst__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_11_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_dst__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_3_en; // @[Decoupled.scala 209:16]
  reg [1:0] ram_msgType [0:1]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_msgType__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_11_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_msgType__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_3_en; // @[Decoupled.scala 209:16]
  reg  enq_ptr_value; // @[Counter.scala 29:33]
  reg  deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = enq_ptr_value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_7 = deq_ptr_value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  wire  _T_10 = ~full; // @[Decoupled.scala 232:19]
  assign ram_addr__T_11_addr = deq_ptr_value;
  assign ram_addr__T_11_data = ram_addr[ram_addr__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_3_data = io_enq_bits_addr;
  assign ram_addr__T_3_addr = enq_ptr_value;
  assign ram_addr__T_3_mask = 1'h1;
  assign ram_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst__T_11_addr = deq_ptr_value;
  assign ram_inst__T_11_data = ram_inst[ram_inst__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst__T_3_data = io_enq_bits_inst;
  assign ram_inst__T_3_addr = enq_ptr_value;
  assign ram_inst__T_3_mask = 1'h1;
  assign ram_inst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_11_addr = deq_ptr_value;
  assign ram_data__T_11_data = ram_data[ram_data__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = enq_ptr_value;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_src__T_11_addr = deq_ptr_value;
  assign ram_src__T_11_data = ram_src[ram_src__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_src__T_3_data = io_enq_bits_src;
  assign ram_src__T_3_addr = enq_ptr_value;
  assign ram_src__T_3_mask = 1'h1;
  assign ram_src__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_dst__T_11_addr = deq_ptr_value;
  assign ram_dst__T_11_data = ram_dst[ram_dst__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_dst__T_3_data = io_enq_bits_dst;
  assign ram_dst__T_3_addr = enq_ptr_value;
  assign ram_dst__T_3_mask = 1'h1;
  assign ram_dst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_msgType__T_11_addr = deq_ptr_value;
  assign ram_msgType__T_11_data = ram_msgType[ram_msgType__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_msgType__T_3_data = io_enq_bits_msgType;
  assign ram_msgType__T_3_addr = enq_ptr_value;
  assign ram_msgType__T_3_mask = 1'h1;
  assign ram_msgType__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | _T_10; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst = ram_inst__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_src = ram_src__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_dst = ram_dst__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_msgType = ram_msgType__T_11_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_inst[initvar] = _RAND_1[7:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_src[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_dst[initvar] = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_msgType[initvar] = _RAND_5[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enq_ptr_value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  deq_ptr_value = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_3_en & ram_addr__T_3_mask) begin
      ram_addr[ram_addr__T_3_addr] <= ram_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst__T_3_en & ram_inst__T_3_mask) begin
      ram_inst[ram_inst__T_3_addr] <= ram_inst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_src__T_3_en & ram_src__T_3_mask) begin
      ram_src[ram_src__T_3_addr] <= ram_src__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_dst__T_3_en & ram_dst__T_3_mask) begin
      ram_dst[ram_dst__T_3_addr] <= ram_dst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_msgType__T_3_en & ram_msgType__T_3_mask) begin
      ram_msgType[ram_msgType__T_3_addr] <= ram_msgType__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 1'h0;
    end else if (do_enq) begin
      enq_ptr_value <= _T_5;
    end
    if (reset) begin
      deq_ptr_value <= 1'h0;
    end else if (do_deq) begin
      deq_ptr_value <= _T_7;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_3(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_inst,
  input  [63:0] io_enq_bits_data,
  input  [2:0]  io_enq_bits_src,
  input  [2:0]  io_enq_bits_dst,
  input  [1:0]  io_enq_bits_msgType,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_inst,
  output [63:0] io_deq_bits_data,
  output [2:0]  io_deq_bits_src,
  output [2:0]  io_deq_bits_dst,
  output [1:0]  io_deq_bits_msgType
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:1]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_11_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [7:0] ram_inst [0:1]; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_11_addr; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_11_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_src [0:1]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_src__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_src__T_11_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_src__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_dst [0:1]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_dst__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_11_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_dst__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_3_en; // @[Decoupled.scala 209:16]
  reg [1:0] ram_msgType [0:1]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_msgType__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_11_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_msgType__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_3_en; // @[Decoupled.scala 209:16]
  reg  enq_ptr_value; // @[Counter.scala 29:33]
  reg  deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = enq_ptr_value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_7 = deq_ptr_value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram_addr__T_11_addr = deq_ptr_value;
  assign ram_addr__T_11_data = ram_addr[ram_addr__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_3_data = io_enq_bits_addr;
  assign ram_addr__T_3_addr = enq_ptr_value;
  assign ram_addr__T_3_mask = 1'h1;
  assign ram_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst__T_11_addr = deq_ptr_value;
  assign ram_inst__T_11_data = ram_inst[ram_inst__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst__T_3_data = io_enq_bits_inst;
  assign ram_inst__T_3_addr = enq_ptr_value;
  assign ram_inst__T_3_mask = 1'h1;
  assign ram_inst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_11_addr = deq_ptr_value;
  assign ram_data__T_11_data = ram_data[ram_data__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = enq_ptr_value;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_src__T_11_addr = deq_ptr_value;
  assign ram_src__T_11_data = ram_src[ram_src__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_src__T_3_data = io_enq_bits_src;
  assign ram_src__T_3_addr = enq_ptr_value;
  assign ram_src__T_3_mask = 1'h1;
  assign ram_src__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_dst__T_11_addr = deq_ptr_value;
  assign ram_dst__T_11_data = ram_dst[ram_dst__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_dst__T_3_data = io_enq_bits_dst;
  assign ram_dst__T_3_addr = enq_ptr_value;
  assign ram_dst__T_3_mask = 1'h1;
  assign ram_dst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_msgType__T_11_addr = deq_ptr_value;
  assign ram_msgType__T_11_data = ram_msgType[ram_msgType__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_msgType__T_3_data = io_enq_bits_msgType;
  assign ram_msgType__T_3_addr = enq_ptr_value;
  assign ram_msgType__T_3_mask = 1'h1;
  assign ram_msgType__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst = ram_inst__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_src = ram_src__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_dst = ram_dst__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_msgType = ram_msgType__T_11_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_inst[initvar] = _RAND_1[7:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_src[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_dst[initvar] = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_msgType[initvar] = _RAND_5[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enq_ptr_value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  deq_ptr_value = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_3_en & ram_addr__T_3_mask) begin
      ram_addr[ram_addr__T_3_addr] <= ram_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst__T_3_en & ram_inst__T_3_mask) begin
      ram_inst[ram_inst__T_3_addr] <= ram_inst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_src__T_3_en & ram_src__T_3_mask) begin
      ram_src[ram_src__T_3_addr] <= ram_src__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_dst__T_3_en & ram_dst__T_3_mask) begin
      ram_dst[ram_dst__T_3_addr] <= ram_dst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_msgType__T_3_en & ram_msgType__T_3_mask) begin
      ram_msgType[ram_msgType__T_3_addr] <= ram_msgType__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 1'h0;
    end else if (do_enq) begin
      enq_ptr_value <= _T_5;
    end
    if (reset) begin
      deq_ptr_value <= 1'h0;
    end else if (do_deq) begin
      deq_ptr_value <= _T_7;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module RRArbiter(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [7:0]  io_in_0_bits_inst,
  input  [63:0] io_in_0_bits_data,
  input  [2:0]  io_in_0_bits_src,
  input  [2:0]  io_in_0_bits_dst,
  input  [1:0]  io_in_0_bits_msgType,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [7:0]  io_in_1_bits_inst,
  input  [63:0] io_in_1_bits_data,
  input  [2:0]  io_in_1_bits_src,
  input  [2:0]  io_in_1_bits_dst,
  input  [1:0]  io_in_1_bits_msgType,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [7:0]  io_out_bits_inst,
  output [63:0] io_out_bits_data,
  output [2:0]  io_out_bits_src,
  output [2:0]  io_out_bits_dst,
  output [1:0]  io_out_bits_msgType,
  output        io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  lastGrant; // @[Reg.scala 15:16]
  wire  grantMask_1 = 1'h1 > lastGrant; // @[Arbiter.scala 67:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbiter.scala 68:75]
  wire  _T_2 = validMask_1 | io_in_0_valid; // @[Arbiter.scala 31:68]
  wire  _T_4 = ~validMask_1; // @[Arbiter.scala 31:78]
  wire  _T_5 = ~_T_2; // @[Arbiter.scala 31:78]
  wire  _T_9 = grantMask_1 | _T_5; // @[Arbiter.scala 72:50]
  wire  _GEN_17 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_4 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_9 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:15]
  assign io_out_bits_inst = io_chosen ? io_in_1_bits_inst : io_in_0_bits_inst; // @[Arbiter.scala 42:15]
  assign io_out_bits_data = io_chosen ? io_in_1_bits_data : io_in_0_bits_data; // @[Arbiter.scala 42:15]
  assign io_out_bits_src = io_chosen ? io_in_1_bits_src : io_in_0_bits_src; // @[Arbiter.scala 42:15]
  assign io_out_bits_dst = io_chosen ? io_in_1_bits_dst : io_in_0_bits_dst; // @[Arbiter.scala 42:15]
  assign io_out_bits_msgType = io_chosen ? io_in_1_bits_msgType : io_in_0_bits_msgType; // @[Arbiter.scala 42:15]
  assign io_chosen = validMask_1 | _GEN_17; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T) begin
      lastGrant <= io_chosen;
    end
  end
endmodule
module Router(
  input         clock,
  input         reset,
  input         io_cacheIn_valid,
  input  [31:0] io_cacheIn_bits_addr,
  input  [7:0]  io_cacheIn_bits_inst,
  input  [63:0] io_cacheIn_bits_data,
  input         io_cacheOut_ready,
  output        io_cacheOut_valid,
  output [31:0] io_cacheOut_bits_addr,
  output [7:0]  io_cacheOut_bits_inst,
  output [63:0] io_cacheOut_bits_data,
  output [1:0]  io_cacheOut_bits_msgType,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [7:0]  io_in_bits_inst,
  input  [63:0] io_in_bits_data,
  input  [2:0]  io_in_bits_src,
  input  [2:0]  io_in_bits_dst,
  input  [1:0]  io_in_bits_msgType,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [7:0]  io_out_bits_inst,
  output [63:0] io_out_bits_data,
  output [2:0]  io_out_bits_src,
  output [2:0]  io_out_bits_dst,
  output [1:0]  io_out_bits_msgType
);
  wire  cache_in_Q_clock; // @[Router.scala 19:26]
  wire  cache_in_Q_reset; // @[Router.scala 19:26]
  wire  cache_in_Q_io_enq_ready; // @[Router.scala 19:26]
  wire  cache_in_Q_io_enq_valid; // @[Router.scala 19:26]
  wire [31:0] cache_in_Q_io_enq_bits_addr; // @[Router.scala 19:26]
  wire [7:0] cache_in_Q_io_enq_bits_inst; // @[Router.scala 19:26]
  wire [63:0] cache_in_Q_io_enq_bits_data; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_enq_bits_src; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_enq_bits_dst; // @[Router.scala 19:26]
  wire [1:0] cache_in_Q_io_enq_bits_msgType; // @[Router.scala 19:26]
  wire  cache_in_Q_io_deq_ready; // @[Router.scala 19:26]
  wire  cache_in_Q_io_deq_valid; // @[Router.scala 19:26]
  wire [31:0] cache_in_Q_io_deq_bits_addr; // @[Router.scala 19:26]
  wire [7:0] cache_in_Q_io_deq_bits_inst; // @[Router.scala 19:26]
  wire [63:0] cache_in_Q_io_deq_bits_data; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_deq_bits_src; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_deq_bits_dst; // @[Router.scala 19:26]
  wire [1:0] cache_in_Q_io_deq_bits_msgType; // @[Router.scala 19:26]
  wire  cache_out_Q_clock; // @[Router.scala 20:27]
  wire  cache_out_Q_reset; // @[Router.scala 20:27]
  wire  cache_out_Q_io_enq_ready; // @[Router.scala 20:27]
  wire  cache_out_Q_io_enq_valid; // @[Router.scala 20:27]
  wire [31:0] cache_out_Q_io_enq_bits_addr; // @[Router.scala 20:27]
  wire [7:0] cache_out_Q_io_enq_bits_inst; // @[Router.scala 20:27]
  wire [63:0] cache_out_Q_io_enq_bits_data; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_enq_bits_src; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_enq_bits_dst; // @[Router.scala 20:27]
  wire [1:0] cache_out_Q_io_enq_bits_msgType; // @[Router.scala 20:27]
  wire  cache_out_Q_io_deq_ready; // @[Router.scala 20:27]
  wire  cache_out_Q_io_deq_valid; // @[Router.scala 20:27]
  wire [31:0] cache_out_Q_io_deq_bits_addr; // @[Router.scala 20:27]
  wire [7:0] cache_out_Q_io_deq_bits_inst; // @[Router.scala 20:27]
  wire [63:0] cache_out_Q_io_deq_bits_data; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_deq_bits_src; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_deq_bits_dst; // @[Router.scala 20:27]
  wire [1:0] cache_out_Q_io_deq_bits_msgType; // @[Router.scala 20:27]
  wire  in_Q_clock; // @[Router.scala 21:20]
  wire  in_Q_reset; // @[Router.scala 21:20]
  wire  in_Q_io_enq_ready; // @[Router.scala 21:20]
  wire  in_Q_io_enq_valid; // @[Router.scala 21:20]
  wire [31:0] in_Q_io_enq_bits_addr; // @[Router.scala 21:20]
  wire [7:0] in_Q_io_enq_bits_inst; // @[Router.scala 21:20]
  wire [63:0] in_Q_io_enq_bits_data; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_enq_bits_src; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_enq_bits_dst; // @[Router.scala 21:20]
  wire [1:0] in_Q_io_enq_bits_msgType; // @[Router.scala 21:20]
  wire  in_Q_io_deq_ready; // @[Router.scala 21:20]
  wire  in_Q_io_deq_valid; // @[Router.scala 21:20]
  wire [31:0] in_Q_io_deq_bits_addr; // @[Router.scala 21:20]
  wire [7:0] in_Q_io_deq_bits_inst; // @[Router.scala 21:20]
  wire [63:0] in_Q_io_deq_bits_data; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_deq_bits_src; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_deq_bits_dst; // @[Router.scala 21:20]
  wire [1:0] in_Q_io_deq_bits_msgType; // @[Router.scala 21:20]
  wire  arbiter_clock; // @[Router.scala 23:23]
  wire  arbiter_io_in_0_ready; // @[Router.scala 23:23]
  wire  arbiter_io_in_0_valid; // @[Router.scala 23:23]
  wire [31:0] arbiter_io_in_0_bits_addr; // @[Router.scala 23:23]
  wire [7:0] arbiter_io_in_0_bits_inst; // @[Router.scala 23:23]
  wire [63:0] arbiter_io_in_0_bits_data; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_0_bits_src; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_0_bits_dst; // @[Router.scala 23:23]
  wire [1:0] arbiter_io_in_0_bits_msgType; // @[Router.scala 23:23]
  wire  arbiter_io_in_1_ready; // @[Router.scala 23:23]
  wire  arbiter_io_in_1_valid; // @[Router.scala 23:23]
  wire [31:0] arbiter_io_in_1_bits_addr; // @[Router.scala 23:23]
  wire [7:0] arbiter_io_in_1_bits_inst; // @[Router.scala 23:23]
  wire [63:0] arbiter_io_in_1_bits_data; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_1_bits_src; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_1_bits_dst; // @[Router.scala 23:23]
  wire [1:0] arbiter_io_in_1_bits_msgType; // @[Router.scala 23:23]
  wire  arbiter_io_out_ready; // @[Router.scala 23:23]
  wire  arbiter_io_out_valid; // @[Router.scala 23:23]
  wire [31:0] arbiter_io_out_bits_addr; // @[Router.scala 23:23]
  wire [7:0] arbiter_io_out_bits_inst; // @[Router.scala 23:23]
  wire [63:0] arbiter_io_out_bits_data; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_out_bits_src; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_out_bits_dst; // @[Router.scala 23:23]
  wire [1:0] arbiter_io_out_bits_msgType; // @[Router.scala 23:23]
  wire  arbiter_io_chosen; // @[Router.scala 23:23]
  wire  _T = in_Q_io_deq_bits_dst == 3'h0; // @[Router.scala 34:74]
  wire  _T_2 = in_Q_io_deq_bits_dst != 3'h0; // @[Router.scala 37:72]
  wire  _T_5 = arbiter_io_in_1_ready & _T_2; // @[Router.scala 38:48]
  wire  _T_7 = cache_out_Q_io_enq_ready & _T; // @[Router.scala 38:113]
  Queue_1 cache_in_Q ( // @[Router.scala 19:26]
    .clock(cache_in_Q_clock),
    .reset(cache_in_Q_reset),
    .io_enq_ready(cache_in_Q_io_enq_ready),
    .io_enq_valid(cache_in_Q_io_enq_valid),
    .io_enq_bits_addr(cache_in_Q_io_enq_bits_addr),
    .io_enq_bits_inst(cache_in_Q_io_enq_bits_inst),
    .io_enq_bits_data(cache_in_Q_io_enq_bits_data),
    .io_enq_bits_src(cache_in_Q_io_enq_bits_src),
    .io_enq_bits_dst(cache_in_Q_io_enq_bits_dst),
    .io_enq_bits_msgType(cache_in_Q_io_enq_bits_msgType),
    .io_deq_ready(cache_in_Q_io_deq_ready),
    .io_deq_valid(cache_in_Q_io_deq_valid),
    .io_deq_bits_addr(cache_in_Q_io_deq_bits_addr),
    .io_deq_bits_inst(cache_in_Q_io_deq_bits_inst),
    .io_deq_bits_data(cache_in_Q_io_deq_bits_data),
    .io_deq_bits_src(cache_in_Q_io_deq_bits_src),
    .io_deq_bits_dst(cache_in_Q_io_deq_bits_dst),
    .io_deq_bits_msgType(cache_in_Q_io_deq_bits_msgType)
  );
  Queue_1 cache_out_Q ( // @[Router.scala 20:27]
    .clock(cache_out_Q_clock),
    .reset(cache_out_Q_reset),
    .io_enq_ready(cache_out_Q_io_enq_ready),
    .io_enq_valid(cache_out_Q_io_enq_valid),
    .io_enq_bits_addr(cache_out_Q_io_enq_bits_addr),
    .io_enq_bits_inst(cache_out_Q_io_enq_bits_inst),
    .io_enq_bits_data(cache_out_Q_io_enq_bits_data),
    .io_enq_bits_src(cache_out_Q_io_enq_bits_src),
    .io_enq_bits_dst(cache_out_Q_io_enq_bits_dst),
    .io_enq_bits_msgType(cache_out_Q_io_enq_bits_msgType),
    .io_deq_ready(cache_out_Q_io_deq_ready),
    .io_deq_valid(cache_out_Q_io_deq_valid),
    .io_deq_bits_addr(cache_out_Q_io_deq_bits_addr),
    .io_deq_bits_inst(cache_out_Q_io_deq_bits_inst),
    .io_deq_bits_data(cache_out_Q_io_deq_bits_data),
    .io_deq_bits_src(cache_out_Q_io_deq_bits_src),
    .io_deq_bits_dst(cache_out_Q_io_deq_bits_dst),
    .io_deq_bits_msgType(cache_out_Q_io_deq_bits_msgType)
  );
  Queue_3 in_Q ( // @[Router.scala 21:20]
    .clock(in_Q_clock),
    .reset(in_Q_reset),
    .io_enq_ready(in_Q_io_enq_ready),
    .io_enq_valid(in_Q_io_enq_valid),
    .io_enq_bits_addr(in_Q_io_enq_bits_addr),
    .io_enq_bits_inst(in_Q_io_enq_bits_inst),
    .io_enq_bits_data(in_Q_io_enq_bits_data),
    .io_enq_bits_src(in_Q_io_enq_bits_src),
    .io_enq_bits_dst(in_Q_io_enq_bits_dst),
    .io_enq_bits_msgType(in_Q_io_enq_bits_msgType),
    .io_deq_ready(in_Q_io_deq_ready),
    .io_deq_valid(in_Q_io_deq_valid),
    .io_deq_bits_addr(in_Q_io_deq_bits_addr),
    .io_deq_bits_inst(in_Q_io_deq_bits_inst),
    .io_deq_bits_data(in_Q_io_deq_bits_data),
    .io_deq_bits_src(in_Q_io_deq_bits_src),
    .io_deq_bits_dst(in_Q_io_deq_bits_dst),
    .io_deq_bits_msgType(in_Q_io_deq_bits_msgType)
  );
  RRArbiter arbiter ( // @[Router.scala 23:23]
    .clock(arbiter_clock),
    .io_in_0_ready(arbiter_io_in_0_ready),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_addr(arbiter_io_in_0_bits_addr),
    .io_in_0_bits_inst(arbiter_io_in_0_bits_inst),
    .io_in_0_bits_data(arbiter_io_in_0_bits_data),
    .io_in_0_bits_src(arbiter_io_in_0_bits_src),
    .io_in_0_bits_dst(arbiter_io_in_0_bits_dst),
    .io_in_0_bits_msgType(arbiter_io_in_0_bits_msgType),
    .io_in_1_ready(arbiter_io_in_1_ready),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_addr(arbiter_io_in_1_bits_addr),
    .io_in_1_bits_inst(arbiter_io_in_1_bits_inst),
    .io_in_1_bits_data(arbiter_io_in_1_bits_data),
    .io_in_1_bits_src(arbiter_io_in_1_bits_src),
    .io_in_1_bits_dst(arbiter_io_in_1_bits_dst),
    .io_in_1_bits_msgType(arbiter_io_in_1_bits_msgType),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_addr(arbiter_io_out_bits_addr),
    .io_out_bits_inst(arbiter_io_out_bits_inst),
    .io_out_bits_data(arbiter_io_out_bits_data),
    .io_out_bits_src(arbiter_io_out_bits_src),
    .io_out_bits_dst(arbiter_io_out_bits_dst),
    .io_out_bits_msgType(arbiter_io_out_bits_msgType),
    .io_chosen(arbiter_io_chosen)
  );
  assign io_cacheOut_valid = cache_out_Q_io_deq_valid; // @[Router.scala 26:15]
  assign io_cacheOut_bits_addr = cache_out_Q_io_deq_bits_addr; // @[Router.scala 26:15]
  assign io_cacheOut_bits_inst = cache_out_Q_io_deq_bits_inst; // @[Router.scala 26:15]
  assign io_cacheOut_bits_data = cache_out_Q_io_deq_bits_data; // @[Router.scala 26:15]
  assign io_cacheOut_bits_msgType = cache_out_Q_io_deq_bits_msgType; // @[Router.scala 26:15]
  assign io_in_ready = in_Q_io_enq_ready; // @[Router.scala 27:15]
  assign io_out_valid = arbiter_io_out_valid; // @[Router.scala 29:10]
  assign io_out_bits_addr = arbiter_io_out_bits_addr; // @[Router.scala 29:10]
  assign io_out_bits_inst = arbiter_io_out_bits_inst; // @[Router.scala 29:10]
  assign io_out_bits_data = arbiter_io_out_bits_data; // @[Router.scala 29:10]
  assign io_out_bits_src = arbiter_io_out_bits_src; // @[Router.scala 29:10]
  assign io_out_bits_dst = arbiter_io_out_bits_dst; // @[Router.scala 29:10]
  assign io_out_bits_msgType = arbiter_io_out_bits_msgType; // @[Router.scala 29:10]
  assign cache_in_Q_clock = clock;
  assign cache_in_Q_reset = reset;
  assign cache_in_Q_io_enq_valid = io_cacheIn_valid; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_addr = io_cacheIn_bits_addr; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_inst = io_cacheIn_bits_inst; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_data = io_cacheIn_bits_data; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_src = 3'h0; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_dst = 3'h1; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_msgType = 2'h0; // @[Router.scala 25:21]
  assign cache_in_Q_io_deq_ready = arbiter_io_in_0_ready; // @[Router.scala 31:20]
  assign cache_out_Q_clock = clock;
  assign cache_out_Q_reset = reset;
  assign cache_out_Q_io_enq_valid = in_Q_io_deq_valid & _T; // @[Router.scala 34:28]
  assign cache_out_Q_io_enq_bits_addr = in_Q_io_deq_bits_addr; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_inst = in_Q_io_deq_bits_inst; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_data = in_Q_io_deq_bits_data; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_src = in_Q_io_deq_bits_src; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_dst = in_Q_io_deq_bits_dst; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_msgType = in_Q_io_deq_bits_msgType; // @[Router.scala 33:27]
  assign cache_out_Q_io_deq_ready = io_cacheOut_ready; // @[Router.scala 26:15]
  assign in_Q_clock = clock;
  assign in_Q_reset = reset;
  assign in_Q_io_enq_valid = io_in_valid; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_addr = io_in_bits_addr; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_inst = io_in_bits_inst; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_data = io_in_bits_data; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_src = io_in_bits_src; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_dst = io_in_bits_dst; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_msgType = io_in_bits_msgType; // @[Router.scala 27:15]
  assign in_Q_io_deq_ready = _T_5 | _T_7; // @[Router.scala 38:21]
  assign arbiter_clock = clock;
  assign arbiter_io_in_0_valid = cache_in_Q_io_deq_valid; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_addr = cache_in_Q_io_deq_bits_addr; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_inst = cache_in_Q_io_deq_bits_inst; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_data = cache_in_Q_io_deq_bits_data; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_src = cache_in_Q_io_deq_bits_src; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_dst = cache_in_Q_io_deq_bits_dst; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_msgType = cache_in_Q_io_deq_bits_msgType; // @[Router.scala 31:20]
  assign arbiter_io_in_1_valid = in_Q_io_deq_valid & _T_2; // @[Router.scala 37:26]
  assign arbiter_io_in_1_bits_addr = in_Q_io_deq_bits_addr; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_inst = in_Q_io_deq_bits_inst; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_data = in_Q_io_deq_bits_data; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_src = in_Q_io_deq_bits_src; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_dst = in_Q_io_deq_bits_dst; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_msgType = in_Q_io_deq_bits_msgType; // @[Router.scala 36:25]
  assign arbiter_io_out_ready = io_out_ready; // @[Router.scala 29:10]
endmodule
module Router_1(
  input         clock,
  input         reset,
  output        io_cacheIn_ready,
  input         io_cacheIn_valid,
  input  [31:0] io_cacheIn_bits_addr,
  input  [63:0] io_cacheIn_bits_data,
  input  [2:0]  io_cacheIn_bits_dst,
  input         io_cacheOut_ready,
  output        io_cacheOut_valid,
  output [31:0] io_cacheOut_bits_addr,
  output [7:0]  io_cacheOut_bits_inst,
  output [63:0] io_cacheOut_bits_data,
  output [2:0]  io_cacheOut_bits_src,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [7:0]  io_in_bits_inst,
  input  [63:0] io_in_bits_data,
  input  [2:0]  io_in_bits_src,
  input  [2:0]  io_in_bits_dst,
  input  [1:0]  io_in_bits_msgType,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [7:0]  io_out_bits_inst,
  output [63:0] io_out_bits_data,
  output [2:0]  io_out_bits_src,
  output [2:0]  io_out_bits_dst,
  output [1:0]  io_out_bits_msgType
);
  wire  cache_in_Q_clock; // @[Router.scala 19:26]
  wire  cache_in_Q_reset; // @[Router.scala 19:26]
  wire  cache_in_Q_io_enq_ready; // @[Router.scala 19:26]
  wire  cache_in_Q_io_enq_valid; // @[Router.scala 19:26]
  wire [31:0] cache_in_Q_io_enq_bits_addr; // @[Router.scala 19:26]
  wire [7:0] cache_in_Q_io_enq_bits_inst; // @[Router.scala 19:26]
  wire [63:0] cache_in_Q_io_enq_bits_data; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_enq_bits_src; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_enq_bits_dst; // @[Router.scala 19:26]
  wire [1:0] cache_in_Q_io_enq_bits_msgType; // @[Router.scala 19:26]
  wire  cache_in_Q_io_deq_ready; // @[Router.scala 19:26]
  wire  cache_in_Q_io_deq_valid; // @[Router.scala 19:26]
  wire [31:0] cache_in_Q_io_deq_bits_addr; // @[Router.scala 19:26]
  wire [7:0] cache_in_Q_io_deq_bits_inst; // @[Router.scala 19:26]
  wire [63:0] cache_in_Q_io_deq_bits_data; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_deq_bits_src; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_deq_bits_dst; // @[Router.scala 19:26]
  wire [1:0] cache_in_Q_io_deq_bits_msgType; // @[Router.scala 19:26]
  wire  cache_out_Q_clock; // @[Router.scala 20:27]
  wire  cache_out_Q_reset; // @[Router.scala 20:27]
  wire  cache_out_Q_io_enq_ready; // @[Router.scala 20:27]
  wire  cache_out_Q_io_enq_valid; // @[Router.scala 20:27]
  wire [31:0] cache_out_Q_io_enq_bits_addr; // @[Router.scala 20:27]
  wire [7:0] cache_out_Q_io_enq_bits_inst; // @[Router.scala 20:27]
  wire [63:0] cache_out_Q_io_enq_bits_data; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_enq_bits_src; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_enq_bits_dst; // @[Router.scala 20:27]
  wire [1:0] cache_out_Q_io_enq_bits_msgType; // @[Router.scala 20:27]
  wire  cache_out_Q_io_deq_ready; // @[Router.scala 20:27]
  wire  cache_out_Q_io_deq_valid; // @[Router.scala 20:27]
  wire [31:0] cache_out_Q_io_deq_bits_addr; // @[Router.scala 20:27]
  wire [7:0] cache_out_Q_io_deq_bits_inst; // @[Router.scala 20:27]
  wire [63:0] cache_out_Q_io_deq_bits_data; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_deq_bits_src; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_deq_bits_dst; // @[Router.scala 20:27]
  wire [1:0] cache_out_Q_io_deq_bits_msgType; // @[Router.scala 20:27]
  wire  in_Q_clock; // @[Router.scala 21:20]
  wire  in_Q_reset; // @[Router.scala 21:20]
  wire  in_Q_io_enq_ready; // @[Router.scala 21:20]
  wire  in_Q_io_enq_valid; // @[Router.scala 21:20]
  wire [31:0] in_Q_io_enq_bits_addr; // @[Router.scala 21:20]
  wire [7:0] in_Q_io_enq_bits_inst; // @[Router.scala 21:20]
  wire [63:0] in_Q_io_enq_bits_data; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_enq_bits_src; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_enq_bits_dst; // @[Router.scala 21:20]
  wire [1:0] in_Q_io_enq_bits_msgType; // @[Router.scala 21:20]
  wire  in_Q_io_deq_ready; // @[Router.scala 21:20]
  wire  in_Q_io_deq_valid; // @[Router.scala 21:20]
  wire [31:0] in_Q_io_deq_bits_addr; // @[Router.scala 21:20]
  wire [7:0] in_Q_io_deq_bits_inst; // @[Router.scala 21:20]
  wire [63:0] in_Q_io_deq_bits_data; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_deq_bits_src; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_deq_bits_dst; // @[Router.scala 21:20]
  wire [1:0] in_Q_io_deq_bits_msgType; // @[Router.scala 21:20]
  wire  arbiter_clock; // @[Router.scala 23:23]
  wire  arbiter_io_in_0_ready; // @[Router.scala 23:23]
  wire  arbiter_io_in_0_valid; // @[Router.scala 23:23]
  wire [31:0] arbiter_io_in_0_bits_addr; // @[Router.scala 23:23]
  wire [7:0] arbiter_io_in_0_bits_inst; // @[Router.scala 23:23]
  wire [63:0] arbiter_io_in_0_bits_data; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_0_bits_src; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_0_bits_dst; // @[Router.scala 23:23]
  wire [1:0] arbiter_io_in_0_bits_msgType; // @[Router.scala 23:23]
  wire  arbiter_io_in_1_ready; // @[Router.scala 23:23]
  wire  arbiter_io_in_1_valid; // @[Router.scala 23:23]
  wire [31:0] arbiter_io_in_1_bits_addr; // @[Router.scala 23:23]
  wire [7:0] arbiter_io_in_1_bits_inst; // @[Router.scala 23:23]
  wire [63:0] arbiter_io_in_1_bits_data; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_1_bits_src; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_1_bits_dst; // @[Router.scala 23:23]
  wire [1:0] arbiter_io_in_1_bits_msgType; // @[Router.scala 23:23]
  wire  arbiter_io_out_ready; // @[Router.scala 23:23]
  wire  arbiter_io_out_valid; // @[Router.scala 23:23]
  wire [31:0] arbiter_io_out_bits_addr; // @[Router.scala 23:23]
  wire [7:0] arbiter_io_out_bits_inst; // @[Router.scala 23:23]
  wire [63:0] arbiter_io_out_bits_data; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_out_bits_src; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_out_bits_dst; // @[Router.scala 23:23]
  wire [1:0] arbiter_io_out_bits_msgType; // @[Router.scala 23:23]
  wire  arbiter_io_chosen; // @[Router.scala 23:23]
  wire  _T = in_Q_io_deq_bits_dst == 3'h1; // @[Router.scala 34:74]
  wire  _T_2 = in_Q_io_deq_bits_dst != 3'h1; // @[Router.scala 37:72]
  wire  _T_5 = arbiter_io_in_1_ready & _T_2; // @[Router.scala 38:48]
  wire  _T_7 = cache_out_Q_io_enq_ready & _T; // @[Router.scala 38:113]
  Queue_1 cache_in_Q ( // @[Router.scala 19:26]
    .clock(cache_in_Q_clock),
    .reset(cache_in_Q_reset),
    .io_enq_ready(cache_in_Q_io_enq_ready),
    .io_enq_valid(cache_in_Q_io_enq_valid),
    .io_enq_bits_addr(cache_in_Q_io_enq_bits_addr),
    .io_enq_bits_inst(cache_in_Q_io_enq_bits_inst),
    .io_enq_bits_data(cache_in_Q_io_enq_bits_data),
    .io_enq_bits_src(cache_in_Q_io_enq_bits_src),
    .io_enq_bits_dst(cache_in_Q_io_enq_bits_dst),
    .io_enq_bits_msgType(cache_in_Q_io_enq_bits_msgType),
    .io_deq_ready(cache_in_Q_io_deq_ready),
    .io_deq_valid(cache_in_Q_io_deq_valid),
    .io_deq_bits_addr(cache_in_Q_io_deq_bits_addr),
    .io_deq_bits_inst(cache_in_Q_io_deq_bits_inst),
    .io_deq_bits_data(cache_in_Q_io_deq_bits_data),
    .io_deq_bits_src(cache_in_Q_io_deq_bits_src),
    .io_deq_bits_dst(cache_in_Q_io_deq_bits_dst),
    .io_deq_bits_msgType(cache_in_Q_io_deq_bits_msgType)
  );
  Queue_1 cache_out_Q ( // @[Router.scala 20:27]
    .clock(cache_out_Q_clock),
    .reset(cache_out_Q_reset),
    .io_enq_ready(cache_out_Q_io_enq_ready),
    .io_enq_valid(cache_out_Q_io_enq_valid),
    .io_enq_bits_addr(cache_out_Q_io_enq_bits_addr),
    .io_enq_bits_inst(cache_out_Q_io_enq_bits_inst),
    .io_enq_bits_data(cache_out_Q_io_enq_bits_data),
    .io_enq_bits_src(cache_out_Q_io_enq_bits_src),
    .io_enq_bits_dst(cache_out_Q_io_enq_bits_dst),
    .io_enq_bits_msgType(cache_out_Q_io_enq_bits_msgType),
    .io_deq_ready(cache_out_Q_io_deq_ready),
    .io_deq_valid(cache_out_Q_io_deq_valid),
    .io_deq_bits_addr(cache_out_Q_io_deq_bits_addr),
    .io_deq_bits_inst(cache_out_Q_io_deq_bits_inst),
    .io_deq_bits_data(cache_out_Q_io_deq_bits_data),
    .io_deq_bits_src(cache_out_Q_io_deq_bits_src),
    .io_deq_bits_dst(cache_out_Q_io_deq_bits_dst),
    .io_deq_bits_msgType(cache_out_Q_io_deq_bits_msgType)
  );
  Queue_3 in_Q ( // @[Router.scala 21:20]
    .clock(in_Q_clock),
    .reset(in_Q_reset),
    .io_enq_ready(in_Q_io_enq_ready),
    .io_enq_valid(in_Q_io_enq_valid),
    .io_enq_bits_addr(in_Q_io_enq_bits_addr),
    .io_enq_bits_inst(in_Q_io_enq_bits_inst),
    .io_enq_bits_data(in_Q_io_enq_bits_data),
    .io_enq_bits_src(in_Q_io_enq_bits_src),
    .io_enq_bits_dst(in_Q_io_enq_bits_dst),
    .io_enq_bits_msgType(in_Q_io_enq_bits_msgType),
    .io_deq_ready(in_Q_io_deq_ready),
    .io_deq_valid(in_Q_io_deq_valid),
    .io_deq_bits_addr(in_Q_io_deq_bits_addr),
    .io_deq_bits_inst(in_Q_io_deq_bits_inst),
    .io_deq_bits_data(in_Q_io_deq_bits_data),
    .io_deq_bits_src(in_Q_io_deq_bits_src),
    .io_deq_bits_dst(in_Q_io_deq_bits_dst),
    .io_deq_bits_msgType(in_Q_io_deq_bits_msgType)
  );
  RRArbiter arbiter ( // @[Router.scala 23:23]
    .clock(arbiter_clock),
    .io_in_0_ready(arbiter_io_in_0_ready),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_addr(arbiter_io_in_0_bits_addr),
    .io_in_0_bits_inst(arbiter_io_in_0_bits_inst),
    .io_in_0_bits_data(arbiter_io_in_0_bits_data),
    .io_in_0_bits_src(arbiter_io_in_0_bits_src),
    .io_in_0_bits_dst(arbiter_io_in_0_bits_dst),
    .io_in_0_bits_msgType(arbiter_io_in_0_bits_msgType),
    .io_in_1_ready(arbiter_io_in_1_ready),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_addr(arbiter_io_in_1_bits_addr),
    .io_in_1_bits_inst(arbiter_io_in_1_bits_inst),
    .io_in_1_bits_data(arbiter_io_in_1_bits_data),
    .io_in_1_bits_src(arbiter_io_in_1_bits_src),
    .io_in_1_bits_dst(arbiter_io_in_1_bits_dst),
    .io_in_1_bits_msgType(arbiter_io_in_1_bits_msgType),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_addr(arbiter_io_out_bits_addr),
    .io_out_bits_inst(arbiter_io_out_bits_inst),
    .io_out_bits_data(arbiter_io_out_bits_data),
    .io_out_bits_src(arbiter_io_out_bits_src),
    .io_out_bits_dst(arbiter_io_out_bits_dst),
    .io_out_bits_msgType(arbiter_io_out_bits_msgType),
    .io_chosen(arbiter_io_chosen)
  );
  assign io_cacheIn_ready = cache_in_Q_io_enq_ready; // @[Router.scala 25:21]
  assign io_cacheOut_valid = cache_out_Q_io_deq_valid; // @[Router.scala 26:15]
  assign io_cacheOut_bits_addr = cache_out_Q_io_deq_bits_addr; // @[Router.scala 26:15]
  assign io_cacheOut_bits_inst = cache_out_Q_io_deq_bits_inst; // @[Router.scala 26:15]
  assign io_cacheOut_bits_data = cache_out_Q_io_deq_bits_data; // @[Router.scala 26:15]
  assign io_cacheOut_bits_src = cache_out_Q_io_deq_bits_src; // @[Router.scala 26:15]
  assign io_in_ready = in_Q_io_enq_ready; // @[Router.scala 27:15]
  assign io_out_valid = arbiter_io_out_valid; // @[Router.scala 29:10]
  assign io_out_bits_addr = arbiter_io_out_bits_addr; // @[Router.scala 29:10]
  assign io_out_bits_inst = arbiter_io_out_bits_inst; // @[Router.scala 29:10]
  assign io_out_bits_data = arbiter_io_out_bits_data; // @[Router.scala 29:10]
  assign io_out_bits_src = arbiter_io_out_bits_src; // @[Router.scala 29:10]
  assign io_out_bits_dst = arbiter_io_out_bits_dst; // @[Router.scala 29:10]
  assign io_out_bits_msgType = arbiter_io_out_bits_msgType; // @[Router.scala 29:10]
  assign cache_in_Q_clock = clock;
  assign cache_in_Q_reset = reset;
  assign cache_in_Q_io_enq_valid = io_cacheIn_valid; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_addr = io_cacheIn_bits_addr; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_inst = 8'h1; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_data = io_cacheIn_bits_data; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_src = 3'h1; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_dst = io_cacheIn_bits_dst; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_msgType = 2'h0; // @[Router.scala 25:21]
  assign cache_in_Q_io_deq_ready = arbiter_io_in_0_ready; // @[Router.scala 31:20]
  assign cache_out_Q_clock = clock;
  assign cache_out_Q_reset = reset;
  assign cache_out_Q_io_enq_valid = in_Q_io_deq_valid & _T; // @[Router.scala 34:28]
  assign cache_out_Q_io_enq_bits_addr = in_Q_io_deq_bits_addr; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_inst = in_Q_io_deq_bits_inst; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_data = in_Q_io_deq_bits_data; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_src = in_Q_io_deq_bits_src; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_dst = in_Q_io_deq_bits_dst; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_msgType = in_Q_io_deq_bits_msgType; // @[Router.scala 33:27]
  assign cache_out_Q_io_deq_ready = io_cacheOut_ready; // @[Router.scala 26:15]
  assign in_Q_clock = clock;
  assign in_Q_reset = reset;
  assign in_Q_io_enq_valid = io_in_valid; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_addr = io_in_bits_addr; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_inst = io_in_bits_inst; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_data = io_in_bits_data; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_src = io_in_bits_src; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_dst = io_in_bits_dst; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_msgType = io_in_bits_msgType; // @[Router.scala 27:15]
  assign in_Q_io_deq_ready = _T_5 | _T_7; // @[Router.scala 38:21]
  assign arbiter_clock = clock;
  assign arbiter_io_in_0_valid = cache_in_Q_io_deq_valid; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_addr = cache_in_Q_io_deq_bits_addr; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_inst = cache_in_Q_io_deq_bits_inst; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_data = cache_in_Q_io_deq_bits_data; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_src = cache_in_Q_io_deq_bits_src; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_dst = cache_in_Q_io_deq_bits_dst; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_msgType = cache_in_Q_io_deq_bits_msgType; // @[Router.scala 31:20]
  assign arbiter_io_in_1_valid = in_Q_io_deq_valid & _T_2; // @[Router.scala 37:26]
  assign arbiter_io_in_1_bits_addr = in_Q_io_deq_bits_addr; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_inst = in_Q_io_deq_bits_inst; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_data = in_Q_io_deq_bits_data; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_src = in_Q_io_deq_bits_src; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_dst = in_Q_io_deq_bits_dst; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_msgType = in_Q_io_deq_bits_msgType; // @[Router.scala 36:25]
  assign arbiter_io_out_ready = io_out_ready; // @[Router.scala 29:10]
endmodule
module bipassLD(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_way,
  output        io_dataMem_in_valid,
  output [31:0] io_dataMem_in_bits_address,
  input  [63:0] io_dataMem_outputValue_0,
  output        io_out_valid,
  output [63:0] io_out_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  set = io_in_bits_addr[0]; // @[Gem5CacheLogic.scala 95:19]
  reg [63:0] dataRead_0; // @[elements.scala 323:27]
  wire [1:0] _GEN_0 = {{1'd0}, set}; // @[elements.scala 327:39]
  wire [2:0] _T_1 = _GEN_0 * 2'h2; // @[elements.scala 327:39]
  wire [2:0] _T_3 = _T_1 + io_in_bits_way; // @[elements.scala 327:49]
  reg  _T_4; // @[elements.scala 331:28]
  assign io_dataMem_in_valid = io_in_valid; // @[elements.scala 325:25]
  assign io_dataMem_in_bits_address = {{29'd0}, _T_3}; // @[elements.scala 327:32]
  assign io_out_valid = _T_4; // @[elements.scala 331:18]
  assign io_out_bits_data = dataRead_0; // @[elements.scala 332:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  dataRead_0 = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  _T_4 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      dataRead_0 <= 64'h0;
    end else begin
      dataRead_0 <= io_dataMem_outputValue_0;
    end
    _T_4 <= io_in_valid;
  end
endmodule
module MemBank(
  input         clock,
  input         io_read_in_valid,
  input  [31:0] io_read_in_bits_address,
  output [63:0] io_read_outputValue_0,
  input         io_write_valid,
  input  [31:0] io_write_bits_address,
  input  [63:0] io_write_bits_inputValue_0
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [63:0] mems_0 [0:3]; // @[BankedMemory.scala 40:8]
  wire [63:0] mems_0__T_1_data; // @[BankedMemory.scala 40:8]
  wire [1:0] mems_0__T_1_addr; // @[BankedMemory.scala 40:8]
  wire [63:0] mems_0__T_5_data; // @[BankedMemory.scala 40:8]
  wire [1:0] mems_0__T_5_addr; // @[BankedMemory.scala 40:8]
  wire  mems_0__T_5_mask; // @[BankedMemory.scala 40:8]
  wire  mems_0__T_5_en; // @[BankedMemory.scala 40:8]
  assign mems_0__T_1_addr = io_read_in_bits_address[1:0];
  assign mems_0__T_1_data = mems_0[mems_0__T_1_addr]; // @[BankedMemory.scala 40:8]
  assign mems_0__T_5_data = io_write_bits_inputValue_0;
  assign mems_0__T_5_addr = io_write_bits_address[1:0];
  assign mems_0__T_5_mask = 1'h1;
  assign mems_0__T_5_en = io_write_valid;
  assign io_read_outputValue_0 = mems_0__T_1_data; // @[BankedMemory.scala 46:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    mems_0[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mems_0__T_5_en & mems_0__T_5_mask) begin
      mems_0[mems_0__T_5_addr] <= mems_0__T_5_data; // @[BankedMemory.scala 40:8]
    end
  end
endmodule
module MemBank_1(
  input         clock,
  input         io_read_in_valid,
  input         io_read_in_bits_address,
  output [30:0] io_read_outputValue_0_tag,
  output [30:0] io_read_outputValue_1_tag,
  input         io_write_valid,
  input  [1:0]  io_write_bits_bank,
  input         io_write_bits_address,
  input  [30:0] io_write_bits_inputValue_0_tag,
  input  [30:0] io_write_bits_inputValue_1_tag
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
  reg [30:0] mems_0_tag [0:1]; // @[BankedMemory.scala 40:8]
  wire [30:0] mems_0_tag__T_data; // @[BankedMemory.scala 40:8]
  wire  mems_0_tag__T_addr; // @[BankedMemory.scala 40:8]
  wire [30:0] mems_0_tag__T_5_data; // @[BankedMemory.scala 40:8]
  wire  mems_0_tag__T_5_addr; // @[BankedMemory.scala 40:8]
  wire  mems_0_tag__T_5_mask; // @[BankedMemory.scala 40:8]
  wire  mems_0_tag__T_5_en; // @[BankedMemory.scala 40:8]
  reg [30:0] mems_1_tag [0:1]; // @[BankedMemory.scala 40:8]
  wire [30:0] mems_1_tag__T_1_data; // @[BankedMemory.scala 40:8]
  wire  mems_1_tag__T_1_addr; // @[BankedMemory.scala 40:8]
  wire [30:0] mems_1_tag__T_9_data; // @[BankedMemory.scala 40:8]
  wire  mems_1_tag__T_9_addr; // @[BankedMemory.scala 40:8]
  wire  mems_1_tag__T_9_mask; // @[BankedMemory.scala 40:8]
  wire  mems_1_tag__T_9_en; // @[BankedMemory.scala 40:8]
  wire  _GEN_17 = io_write_bits_bank[0] ? 1'h0 : io_write_bits_bank[1]; // @[BankedMemory.scala 57:82]
  assign mems_0_tag__T_addr = io_read_in_bits_address;
  assign mems_0_tag__T_data = mems_0_tag[mems_0_tag__T_addr]; // @[BankedMemory.scala 40:8]
  assign mems_0_tag__T_5_data = io_write_bits_inputValue_0_tag;
  assign mems_0_tag__T_5_addr = io_write_bits_address;
  assign mems_0_tag__T_5_mask = 1'h1;
  assign mems_0_tag__T_5_en = io_write_valid & io_write_bits_bank[0];
  assign mems_1_tag__T_1_addr = io_read_in_bits_address;
  assign mems_1_tag__T_1_data = mems_1_tag[mems_1_tag__T_1_addr]; // @[BankedMemory.scala 40:8]
  assign mems_1_tag__T_9_data = io_write_bits_inputValue_1_tag;
  assign mems_1_tag__T_9_addr = io_write_bits_address;
  assign mems_1_tag__T_9_mask = 1'h1;
  assign mems_1_tag__T_9_en = io_write_valid & _GEN_17;
  assign io_read_outputValue_0_tag = mems_0_tag__T_data; // @[BankedMemory.scala 46:42]
  assign io_read_outputValue_1_tag = mems_1_tag__T_1_data; // @[BankedMemory.scala 46:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    mems_0_tag[initvar] = _RAND_0[30:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    mems_1_tag[initvar] = _RAND_1[30:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mems_0_tag__T_5_en & mems_0_tag__T_5_mask) begin
      mems_0_tag[mems_0_tag__T_5_addr] <= mems_0_tag__T_5_data; // @[BankedMemory.scala 40:8]
    end
    if(mems_1_tag__T_9_en & mems_1_tag__T_9_mask) begin
      mems_1_tag[mems_1_tag__T_9_addr] <= mems_1_tag__T_9_data; // @[BankedMemory.scala 40:8]
    end
  end
endmodule
module Decoder(
  input  [27:0] io_inAction,
  output        io_outSignals_0,
  output        io_outSignals_1,
  output        io_outSignals_2,
  output        io_outSignals_3,
  output        io_outSignals_4,
  output        io_outSignals_5,
  output        io_outSignals_6,
  output        io_outSignals_7,
  output        io_outSignals_8
);
  assign io_outSignals_0 = io_inAction[0]; // @[elements.scala 21:19]
  assign io_outSignals_1 = io_inAction[1]; // @[elements.scala 21:19]
  assign io_outSignals_2 = io_inAction[2]; // @[elements.scala 21:19]
  assign io_outSignals_3 = io_inAction[3]; // @[elements.scala 21:19]
  assign io_outSignals_4 = io_inAction[4]; // @[elements.scala 21:19]
  assign io_outSignals_5 = io_inAction[5]; // @[elements.scala 21:19]
  assign io_outSignals_6 = io_inAction[6]; // @[elements.scala 21:19]
  assign io_outSignals_7 = io_inAction[7]; // @[elements.scala 21:19]
  assign io_outSignals_8 = io_inAction[8]; // @[elements.scala 21:19]
endmodule
module FindEmptyLine(
  input   io_data_0,
  input   io_data_1,
  output  io_value_valid
);
  wire  _T = ~io_data_0; // @[elements.scala 74:53]
  wire  _T_1 = ~io_data_1; // @[elements.scala 74:53]
  assign io_value_valid = _T | _T_1; // @[elements.scala 68:20 elements.scala 76:32 elements.scala 76:32]
endmodule
module Find(
  input  [30:0] io_key_tag,
  input  [30:0] io_data_0_tag,
  input  [30:0] io_data_1_tag,
  input         io_valid_0,
  input         io_valid_1,
  output        io_value_valid,
  output [31:0] io_value_bits
);
  wire  _T = io_data_0_tag == io_key_tag; // @[elements.scala 35:54]
  wire  _T_1 = io_data_1_tag == io_key_tag; // @[elements.scala 35:54]
  wire [1:0] bitmap = {_T_1,_T}; // @[Cat.scala 29:58]
  wire [1:0] _T_3 = {io_valid_1,io_valid_0}; // @[elements.scala 36:46]
  wire [1:0] _T_4 = bitmap & _T_3; // @[elements.scala 36:29]
  assign io_value_valid = _T_4 != 2'h0; // @[elements.scala 39:20]
  assign io_value_bits = {{31'd0}, _T_4[1]}; // @[elements.scala 38:19]
endmodule
module Gem5CacheLogic(
  input         clock,
  input         reset,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [27:0] io_cpu_req_bits_command,
  input  [1:0]  io_cpu_req_bits_way,
  input  [1:0]  io_cpu_req_bits_replaceWay,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_iswrite,
  output [1:0]  io_cpu_resp_bits_way,
  output        io_metaMem_write_valid,
  output [1:0]  io_metaMem_write_bits_bank,
  output        io_metaMem_write_bits_address,
  output [30:0] io_metaMem_write_bits_inputValue_0_tag,
  output [30:0] io_metaMem_write_bits_inputValue_1_tag,
  output        io_validTagBits_write_valid,
  output [63:0] io_validTagBits_write_bits_addr,
  output        io_validTagBits_write_bits_value,
  output        io_validTagBits_read_in_valid,
  output [63:0] io_validTagBits_read_in_bits_addr,
  input         io_validTagBits_read_out_0,
  input         io_validTagBits_read_out_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [27:0] decoder_io_inAction; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_7; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_8; // @[Gem5CacheLogic.scala 188:23]
  wire  emptyLine_io_data_0; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_data_1; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 359:25]
  wire [30:0] tagFinder_io_key_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_0_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_1_tag; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_0; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_1; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_value_valid; // @[Gem5CacheLogic.scala 362:25]
  wire [31:0] tagFinder_io_value_bits; // @[Gem5CacheLogic.scala 362:25]
  reg [31:0] addr_reg; // @[Gem5CacheLogic.scala 202:25]
  reg [27:0] cpu_command; // @[Gem5CacheLogic.scala 205:28]
  reg [30:0] tag; // @[Gem5CacheLogic.scala 207:20]
  reg  set; // @[Gem5CacheLogic.scala 208:20]
  reg [2:0] wayInput; // @[Gem5CacheLogic.scala 209:25]
  reg [2:0] replaceWayInput; // @[Gem5CacheLogic.scala 210:32]
  wire  _T_3 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_47 = {{1'd0}, set}; // @[Gem5CacheLogic.scala 289:41]
  wire [2:0] _T_6 = _GEN_47 * 2'h2; // @[Gem5CacheLogic.scala 289:41]
  wire  signals_2 = decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  wayInvalid = wayInput == 3'h2; // @[Gem5CacheLogic.scala 351:27]
  wire  _T_28 = ~wayInvalid; // @[Gem5CacheLogic.scala 378:14]
  wire [2:0] _GEN_15 = _T_28 ? wayInput : 3'h2; // @[Gem5CacheLogic.scala 378:26]
  wire [2:0] way = signals_2 ? replaceWayInput : _GEN_15; // @[Gem5CacheLogic.scala 376:23]
  wire [2:0] _T_8 = _T_6 + way; // @[Gem5CacheLogic.scala 289:51]
  wire  signals_1 = decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_0 = decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_23 = signals_1 & signals_0; // @[Gem5CacheLogic.scala 367:37]
  wire  _T_24 = signals_2 | _T_23; // @[Gem5CacheLogic.scala 367:21]
  wire [2:0] _GEN_14 = _T_24 ? _T_6 : 3'h0; // @[Gem5CacheLogic.scala 367:53]
  wire [7:0] _T_29 = 8'h1 << way; // @[Gem5CacheLogic.scala 338:34]
  wire  signals_4 = decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_3 = decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire [31:0] _T_47 = tagFinder_io_value_valid ? tagFinder_io_value_bits : 32'h2; // @[Gem5CacheLogic.scala 424:25]
  wire [2:0] _GEN_41 = signals_2 ? way : 3'h2; // @[Gem5CacheLogic.scala 425:28]
  wire [31:0] _GEN_43 = _T_23 ? _T_47 : {{29'd0}, _GEN_41}; // @[Gem5CacheLogic.scala 423:39]
  wire  signals_5 = decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_6 = decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_52 = ~signals_6; // @[Gem5CacheLogic.scala 446:50]
  reg  _T_54; // @[Gem5CacheLogic.scala 455:38]
  reg  _T_57; // @[Gem5CacheLogic.scala 456:81]
  wire  _T_59 = ~emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 460:26]
  wire  _T_60 = signals_2 & _T_59; // @[Gem5CacheLogic.scala 460:23]
  wire  _T_62 = ~reset; // @[Gem5CacheLogic.scala 461:13]
  wire [2:0] targetWayWire = _GEN_43[2:0]; // @[Gem5CacheLogic.scala 424:19 Gem5CacheLogic.scala 426:19]
  Decoder decoder ( // @[Gem5CacheLogic.scala 188:23]
    .io_inAction(decoder_io_inAction),
    .io_outSignals_0(decoder_io_outSignals_0),
    .io_outSignals_1(decoder_io_outSignals_1),
    .io_outSignals_2(decoder_io_outSignals_2),
    .io_outSignals_3(decoder_io_outSignals_3),
    .io_outSignals_4(decoder_io_outSignals_4),
    .io_outSignals_5(decoder_io_outSignals_5),
    .io_outSignals_6(decoder_io_outSignals_6),
    .io_outSignals_7(decoder_io_outSignals_7),
    .io_outSignals_8(decoder_io_outSignals_8)
  );
  FindEmptyLine emptyLine ( // @[Gem5CacheLogic.scala 359:25]
    .io_data_0(emptyLine_io_data_0),
    .io_data_1(emptyLine_io_data_1),
    .io_value_valid(emptyLine_io_value_valid)
  );
  Find tagFinder ( // @[Gem5CacheLogic.scala 362:25]
    .io_key_tag(tagFinder_io_key_tag),
    .io_data_0_tag(tagFinder_io_data_0_tag),
    .io_data_1_tag(tagFinder_io_data_1_tag),
    .io_valid_0(tagFinder_io_valid_0),
    .io_valid_1(tagFinder_io_valid_1),
    .io_value_valid(tagFinder_io_value_valid),
    .io_value_bits(tagFinder_io_value_bits)
  );
  assign io_cpu_req_ready = 1'h1; // @[Gem5CacheLogic.scala 302:20]
  assign io_cpu_resp_valid = _T_24 | _T_57; // @[Gem5CacheLogic.scala 456:24]
  assign io_cpu_resp_bits_iswrite = _T_54; // @[Gem5CacheLogic.scala 455:28]
  assign io_cpu_resp_bits_way = targetWayWire[1:0]; // @[Gem5CacheLogic.scala 453:24]
  assign io_metaMem_write_valid = signals_3 ? 1'h0 : signals_4; // @[Gem5CacheLogic.scala 346:26 Gem5CacheLogic.scala 330:19]
  assign io_metaMem_write_bits_bank = _T_29[1:0]; // @[Gem5CacheLogic.scala 338:27]
  assign io_metaMem_write_bits_address = set; // @[Gem5CacheLogic.scala 339:30]
  assign io_metaMem_write_bits_inputValue_0_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_metaMem_write_bits_inputValue_1_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_validTagBits_write_valid = signals_5 | signals_6; // @[Gem5CacheLogic.scala 445:31]
  assign io_validTagBits_write_bits_addr = {{61'd0}, _T_8}; // @[Gem5CacheLogic.scala 444:35]
  assign io_validTagBits_write_bits_value = signals_5 | _T_52; // @[Gem5CacheLogic.scala 446:36]
  assign io_validTagBits_read_in_valid = signals_2 | _T_23; // @[Gem5CacheLogic.scala 373:33]
  assign io_validTagBits_read_in_bits_addr = {{61'd0}, _GEN_14}; // @[Gem5CacheLogic.scala 368:39 Gem5CacheLogic.scala 370:39]
  assign decoder_io_inAction = cpu_command; // @[Gem5CacheLogic.scala 298:23]
  assign emptyLine_io_data_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 360:21]
  assign emptyLine_io_data_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 360:21]
  assign tagFinder_io_key_tag = tag; // @[Gem5CacheLogic.scala 363:20]
  assign tagFinder_io_data_0_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_data_1_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_valid_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 365:22]
  assign tagFinder_io_valid_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 365:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cpu_command = _RAND_1[27:0];
  _RAND_2 = {1{`RANDOM}};
  tag = _RAND_2[30:0];
  _RAND_3 = {1{`RANDOM}};
  set = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wayInput = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  replaceWayInput = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _T_54 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_57 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr_reg <= 32'h0;
    end else if (_T_3) begin
      addr_reg <= io_cpu_req_bits_addr;
    end
    if (reset) begin
      cpu_command <= 28'h0;
    end else if (_T_3) begin
      cpu_command <= io_cpu_req_bits_command;
    end
    if (reset) begin
      tag <= 31'h0;
    end else if (_T_3) begin
      tag <= io_cpu_req_bits_addr[31:1];
    end
    if (reset) begin
      set <= 1'h0;
    end else if (_T_3) begin
      set <= io_cpu_req_bits_addr[0];
    end
    if (reset) begin
      wayInput <= 3'h2;
    end else if (_T_3) begin
      wayInput <= {{1'd0}, io_cpu_req_bits_way};
    end
    if (reset) begin
      replaceWayInput <= 3'h2;
    end else if (_T_3) begin
      replaceWayInput <= {{1'd0}, io_cpu_req_bits_replaceWay};
    end
    _T_54 <= decoder_io_outSignals_8;
    _T_57 <= decoder_io_outSignals_8;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_60 & _T_62) begin
          $fwrite(32'h80000002,"Replacement in Set: %d, Way: %d, Addr: %d\n",set,way,addr_reg); // @[Gem5CacheLogic.scala 461:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Gem5CacheLogic_1(
  input         clock,
  input         reset,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [27:0] io_cpu_req_bits_command,
  input  [1:0]  io_cpu_req_bits_way,
  input  [1:0]  io_cpu_req_bits_replaceWay,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_iswrite,
  output [1:0]  io_cpu_resp_bits_way,
  output        io_metaMem_write_valid,
  output [1:0]  io_metaMem_write_bits_bank,
  output        io_metaMem_write_bits_address,
  output [30:0] io_metaMem_write_bits_inputValue_0_tag,
  output [30:0] io_metaMem_write_bits_inputValue_1_tag,
  output        io_validTagBits_write_valid,
  output [63:0] io_validTagBits_write_bits_addr,
  output        io_validTagBits_write_bits_value,
  output        io_validTagBits_read_in_valid,
  output [63:0] io_validTagBits_read_in_bits_addr,
  input         io_validTagBits_read_out_0,
  input         io_validTagBits_read_out_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [27:0] decoder_io_inAction; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_7; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_8; // @[Gem5CacheLogic.scala 188:23]
  wire  emptyLine_io_data_0; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_data_1; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 359:25]
  wire [30:0] tagFinder_io_key_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_0_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_1_tag; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_0; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_1; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_value_valid; // @[Gem5CacheLogic.scala 362:25]
  wire [31:0] tagFinder_io_value_bits; // @[Gem5CacheLogic.scala 362:25]
  reg [31:0] addr_reg; // @[Gem5CacheLogic.scala 202:25]
  reg [27:0] cpu_command; // @[Gem5CacheLogic.scala 205:28]
  reg [30:0] tag; // @[Gem5CacheLogic.scala 207:20]
  reg  set; // @[Gem5CacheLogic.scala 208:20]
  reg [2:0] wayInput; // @[Gem5CacheLogic.scala 209:25]
  reg [2:0] replaceWayInput; // @[Gem5CacheLogic.scala 210:32]
  wire  _T_3 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_47 = {{1'd0}, set}; // @[Gem5CacheLogic.scala 289:41]
  wire [2:0] _T_6 = _GEN_47 * 2'h2; // @[Gem5CacheLogic.scala 289:41]
  wire  signals_2 = decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  wayInvalid = wayInput == 3'h2; // @[Gem5CacheLogic.scala 351:27]
  wire  _T_28 = ~wayInvalid; // @[Gem5CacheLogic.scala 378:14]
  wire [2:0] _GEN_15 = _T_28 ? wayInput : 3'h2; // @[Gem5CacheLogic.scala 378:26]
  wire [2:0] way = signals_2 ? replaceWayInput : _GEN_15; // @[Gem5CacheLogic.scala 376:23]
  wire [2:0] _T_8 = _T_6 + way; // @[Gem5CacheLogic.scala 289:51]
  wire  signals_1 = decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_0 = decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_23 = signals_1 & signals_0; // @[Gem5CacheLogic.scala 367:37]
  wire  _T_24 = signals_2 | _T_23; // @[Gem5CacheLogic.scala 367:21]
  wire [2:0] _GEN_14 = _T_24 ? _T_6 : 3'h0; // @[Gem5CacheLogic.scala 367:53]
  wire [7:0] _T_29 = 8'h1 << way; // @[Gem5CacheLogic.scala 338:34]
  wire  signals_4 = decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_3 = decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire [31:0] _T_47 = tagFinder_io_value_valid ? tagFinder_io_value_bits : 32'h2; // @[Gem5CacheLogic.scala 424:25]
  wire [2:0] _GEN_41 = signals_2 ? way : 3'h2; // @[Gem5CacheLogic.scala 425:28]
  wire [31:0] _GEN_43 = _T_23 ? _T_47 : {{29'd0}, _GEN_41}; // @[Gem5CacheLogic.scala 423:39]
  wire  signals_5 = decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_6 = decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_52 = ~signals_6; // @[Gem5CacheLogic.scala 446:50]
  reg  _T_54; // @[Gem5CacheLogic.scala 455:38]
  reg  _T_57; // @[Gem5CacheLogic.scala 456:81]
  wire  _T_59 = ~emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 460:26]
  wire  _T_60 = signals_2 & _T_59; // @[Gem5CacheLogic.scala 460:23]
  wire  _T_62 = ~reset; // @[Gem5CacheLogic.scala 461:13]
  wire [2:0] targetWayWire = _GEN_43[2:0]; // @[Gem5CacheLogic.scala 424:19 Gem5CacheLogic.scala 426:19]
  Decoder decoder ( // @[Gem5CacheLogic.scala 188:23]
    .io_inAction(decoder_io_inAction),
    .io_outSignals_0(decoder_io_outSignals_0),
    .io_outSignals_1(decoder_io_outSignals_1),
    .io_outSignals_2(decoder_io_outSignals_2),
    .io_outSignals_3(decoder_io_outSignals_3),
    .io_outSignals_4(decoder_io_outSignals_4),
    .io_outSignals_5(decoder_io_outSignals_5),
    .io_outSignals_6(decoder_io_outSignals_6),
    .io_outSignals_7(decoder_io_outSignals_7),
    .io_outSignals_8(decoder_io_outSignals_8)
  );
  FindEmptyLine emptyLine ( // @[Gem5CacheLogic.scala 359:25]
    .io_data_0(emptyLine_io_data_0),
    .io_data_1(emptyLine_io_data_1),
    .io_value_valid(emptyLine_io_value_valid)
  );
  Find tagFinder ( // @[Gem5CacheLogic.scala 362:25]
    .io_key_tag(tagFinder_io_key_tag),
    .io_data_0_tag(tagFinder_io_data_0_tag),
    .io_data_1_tag(tagFinder_io_data_1_tag),
    .io_valid_0(tagFinder_io_valid_0),
    .io_valid_1(tagFinder_io_valid_1),
    .io_value_valid(tagFinder_io_value_valid),
    .io_value_bits(tagFinder_io_value_bits)
  );
  assign io_cpu_req_ready = 1'h1; // @[Gem5CacheLogic.scala 302:20]
  assign io_cpu_resp_valid = _T_24 | _T_57; // @[Gem5CacheLogic.scala 456:24]
  assign io_cpu_resp_bits_iswrite = _T_54; // @[Gem5CacheLogic.scala 455:28]
  assign io_cpu_resp_bits_way = targetWayWire[1:0]; // @[Gem5CacheLogic.scala 453:24]
  assign io_metaMem_write_valid = signals_3 ? 1'h0 : signals_4; // @[Gem5CacheLogic.scala 346:26 Gem5CacheLogic.scala 330:19]
  assign io_metaMem_write_bits_bank = _T_29[1:0]; // @[Gem5CacheLogic.scala 338:27]
  assign io_metaMem_write_bits_address = set; // @[Gem5CacheLogic.scala 339:30]
  assign io_metaMem_write_bits_inputValue_0_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_metaMem_write_bits_inputValue_1_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_validTagBits_write_valid = signals_5 | signals_6; // @[Gem5CacheLogic.scala 445:31]
  assign io_validTagBits_write_bits_addr = {{61'd0}, _T_8}; // @[Gem5CacheLogic.scala 444:35]
  assign io_validTagBits_write_bits_value = signals_5 | _T_52; // @[Gem5CacheLogic.scala 446:36]
  assign io_validTagBits_read_in_valid = signals_2 | _T_23; // @[Gem5CacheLogic.scala 373:33]
  assign io_validTagBits_read_in_bits_addr = {{61'd0}, _GEN_14}; // @[Gem5CacheLogic.scala 368:39 Gem5CacheLogic.scala 370:39]
  assign decoder_io_inAction = cpu_command; // @[Gem5CacheLogic.scala 298:23]
  assign emptyLine_io_data_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 360:21]
  assign emptyLine_io_data_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 360:21]
  assign tagFinder_io_key_tag = tag; // @[Gem5CacheLogic.scala 363:20]
  assign tagFinder_io_data_0_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_data_1_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_valid_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 365:22]
  assign tagFinder_io_valid_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 365:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cpu_command = _RAND_1[27:0];
  _RAND_2 = {1{`RANDOM}};
  tag = _RAND_2[30:0];
  _RAND_3 = {1{`RANDOM}};
  set = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wayInput = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  replaceWayInput = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _T_54 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_57 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr_reg <= 32'h0;
    end else if (_T_3) begin
      addr_reg <= io_cpu_req_bits_addr;
    end
    if (reset) begin
      cpu_command <= 28'h0;
    end else if (_T_3) begin
      cpu_command <= io_cpu_req_bits_command;
    end
    if (reset) begin
      tag <= 31'h0;
    end else if (_T_3) begin
      tag <= io_cpu_req_bits_addr[31:1];
    end
    if (reset) begin
      set <= 1'h0;
    end else if (_T_3) begin
      set <= io_cpu_req_bits_addr[0];
    end
    if (reset) begin
      wayInput <= 3'h2;
    end else if (_T_3) begin
      wayInput <= {{1'd0}, io_cpu_req_bits_way};
    end
    if (reset) begin
      replaceWayInput <= 3'h2;
    end else if (_T_3) begin
      replaceWayInput <= {{1'd0}, io_cpu_req_bits_replaceWay};
    end
    _T_54 <= decoder_io_outSignals_8;
    _T_57 <= decoder_io_outSignals_8;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_60 & _T_62) begin
          $fwrite(32'h80000002,"Replacement in Set: %d, Way: %d, Addr: %d\n",set,way,addr_reg); // @[Gem5CacheLogic.scala 461:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Gem5CacheLogic_2(
  input         clock,
  input         reset,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [27:0] io_cpu_req_bits_command,
  input  [1:0]  io_cpu_req_bits_way,
  input  [1:0]  io_cpu_req_bits_replaceWay,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_iswrite,
  output [1:0]  io_cpu_resp_bits_way,
  output        io_metaMem_write_valid,
  output [1:0]  io_metaMem_write_bits_bank,
  output        io_metaMem_write_bits_address,
  output [30:0] io_metaMem_write_bits_inputValue_0_tag,
  output [30:0] io_metaMem_write_bits_inputValue_1_tag,
  output        io_validTagBits_write_valid,
  output [63:0] io_validTagBits_write_bits_addr,
  output        io_validTagBits_write_bits_value,
  output        io_validTagBits_read_in_valid,
  output [63:0] io_validTagBits_read_in_bits_addr,
  input         io_validTagBits_read_out_0,
  input         io_validTagBits_read_out_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [27:0] decoder_io_inAction; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_7; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_8; // @[Gem5CacheLogic.scala 188:23]
  wire  emptyLine_io_data_0; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_data_1; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 359:25]
  wire [30:0] tagFinder_io_key_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_0_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_1_tag; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_0; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_1; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_value_valid; // @[Gem5CacheLogic.scala 362:25]
  wire [31:0] tagFinder_io_value_bits; // @[Gem5CacheLogic.scala 362:25]
  reg [31:0] addr_reg; // @[Gem5CacheLogic.scala 202:25]
  reg [27:0] cpu_command; // @[Gem5CacheLogic.scala 205:28]
  reg [30:0] tag; // @[Gem5CacheLogic.scala 207:20]
  reg  set; // @[Gem5CacheLogic.scala 208:20]
  reg [2:0] wayInput; // @[Gem5CacheLogic.scala 209:25]
  reg [2:0] replaceWayInput; // @[Gem5CacheLogic.scala 210:32]
  wire  _T_3 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_47 = {{1'd0}, set}; // @[Gem5CacheLogic.scala 289:41]
  wire [2:0] _T_6 = _GEN_47 * 2'h2; // @[Gem5CacheLogic.scala 289:41]
  wire  signals_2 = decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  wayInvalid = wayInput == 3'h2; // @[Gem5CacheLogic.scala 351:27]
  wire  _T_28 = ~wayInvalid; // @[Gem5CacheLogic.scala 378:14]
  wire [2:0] _GEN_15 = _T_28 ? wayInput : 3'h2; // @[Gem5CacheLogic.scala 378:26]
  wire [2:0] way = signals_2 ? replaceWayInput : _GEN_15; // @[Gem5CacheLogic.scala 376:23]
  wire [2:0] _T_8 = _T_6 + way; // @[Gem5CacheLogic.scala 289:51]
  wire  signals_1 = decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_0 = decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_23 = signals_1 & signals_0; // @[Gem5CacheLogic.scala 367:37]
  wire  _T_24 = signals_2 | _T_23; // @[Gem5CacheLogic.scala 367:21]
  wire [2:0] _GEN_14 = _T_24 ? _T_6 : 3'h0; // @[Gem5CacheLogic.scala 367:53]
  wire [7:0] _T_29 = 8'h1 << way; // @[Gem5CacheLogic.scala 338:34]
  wire  signals_4 = decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_3 = decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire [31:0] _T_47 = tagFinder_io_value_valid ? tagFinder_io_value_bits : 32'h2; // @[Gem5CacheLogic.scala 424:25]
  wire [2:0] _GEN_41 = signals_2 ? way : 3'h2; // @[Gem5CacheLogic.scala 425:28]
  wire [31:0] _GEN_43 = _T_23 ? _T_47 : {{29'd0}, _GEN_41}; // @[Gem5CacheLogic.scala 423:39]
  wire  signals_5 = decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_6 = decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_52 = ~signals_6; // @[Gem5CacheLogic.scala 446:50]
  reg  _T_54; // @[Gem5CacheLogic.scala 455:38]
  reg  _T_57; // @[Gem5CacheLogic.scala 456:81]
  wire  _T_59 = ~emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 460:26]
  wire  _T_60 = signals_2 & _T_59; // @[Gem5CacheLogic.scala 460:23]
  wire  _T_62 = ~reset; // @[Gem5CacheLogic.scala 461:13]
  wire [2:0] targetWayWire = _GEN_43[2:0]; // @[Gem5CacheLogic.scala 424:19 Gem5CacheLogic.scala 426:19]
  Decoder decoder ( // @[Gem5CacheLogic.scala 188:23]
    .io_inAction(decoder_io_inAction),
    .io_outSignals_0(decoder_io_outSignals_0),
    .io_outSignals_1(decoder_io_outSignals_1),
    .io_outSignals_2(decoder_io_outSignals_2),
    .io_outSignals_3(decoder_io_outSignals_3),
    .io_outSignals_4(decoder_io_outSignals_4),
    .io_outSignals_5(decoder_io_outSignals_5),
    .io_outSignals_6(decoder_io_outSignals_6),
    .io_outSignals_7(decoder_io_outSignals_7),
    .io_outSignals_8(decoder_io_outSignals_8)
  );
  FindEmptyLine emptyLine ( // @[Gem5CacheLogic.scala 359:25]
    .io_data_0(emptyLine_io_data_0),
    .io_data_1(emptyLine_io_data_1),
    .io_value_valid(emptyLine_io_value_valid)
  );
  Find tagFinder ( // @[Gem5CacheLogic.scala 362:25]
    .io_key_tag(tagFinder_io_key_tag),
    .io_data_0_tag(tagFinder_io_data_0_tag),
    .io_data_1_tag(tagFinder_io_data_1_tag),
    .io_valid_0(tagFinder_io_valid_0),
    .io_valid_1(tagFinder_io_valid_1),
    .io_value_valid(tagFinder_io_value_valid),
    .io_value_bits(tagFinder_io_value_bits)
  );
  assign io_cpu_req_ready = 1'h1; // @[Gem5CacheLogic.scala 302:20]
  assign io_cpu_resp_valid = _T_24 | _T_57; // @[Gem5CacheLogic.scala 456:24]
  assign io_cpu_resp_bits_iswrite = _T_54; // @[Gem5CacheLogic.scala 455:28]
  assign io_cpu_resp_bits_way = targetWayWire[1:0]; // @[Gem5CacheLogic.scala 453:24]
  assign io_metaMem_write_valid = signals_3 ? 1'h0 : signals_4; // @[Gem5CacheLogic.scala 346:26 Gem5CacheLogic.scala 330:19]
  assign io_metaMem_write_bits_bank = _T_29[1:0]; // @[Gem5CacheLogic.scala 338:27]
  assign io_metaMem_write_bits_address = set; // @[Gem5CacheLogic.scala 339:30]
  assign io_metaMem_write_bits_inputValue_0_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_metaMem_write_bits_inputValue_1_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_validTagBits_write_valid = signals_5 | signals_6; // @[Gem5CacheLogic.scala 445:31]
  assign io_validTagBits_write_bits_addr = {{61'd0}, _T_8}; // @[Gem5CacheLogic.scala 444:35]
  assign io_validTagBits_write_bits_value = signals_5 | _T_52; // @[Gem5CacheLogic.scala 446:36]
  assign io_validTagBits_read_in_valid = signals_2 | _T_23; // @[Gem5CacheLogic.scala 373:33]
  assign io_validTagBits_read_in_bits_addr = {{61'd0}, _GEN_14}; // @[Gem5CacheLogic.scala 368:39 Gem5CacheLogic.scala 370:39]
  assign decoder_io_inAction = cpu_command; // @[Gem5CacheLogic.scala 298:23]
  assign emptyLine_io_data_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 360:21]
  assign emptyLine_io_data_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 360:21]
  assign tagFinder_io_key_tag = tag; // @[Gem5CacheLogic.scala 363:20]
  assign tagFinder_io_data_0_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_data_1_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_valid_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 365:22]
  assign tagFinder_io_valid_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 365:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cpu_command = _RAND_1[27:0];
  _RAND_2 = {1{`RANDOM}};
  tag = _RAND_2[30:0];
  _RAND_3 = {1{`RANDOM}};
  set = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wayInput = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  replaceWayInput = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _T_54 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_57 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr_reg <= 32'h0;
    end else if (_T_3) begin
      addr_reg <= io_cpu_req_bits_addr;
    end
    if (reset) begin
      cpu_command <= 28'h0;
    end else if (_T_3) begin
      cpu_command <= io_cpu_req_bits_command;
    end
    if (reset) begin
      tag <= 31'h0;
    end else if (_T_3) begin
      tag <= io_cpu_req_bits_addr[31:1];
    end
    if (reset) begin
      set <= 1'h0;
    end else if (_T_3) begin
      set <= io_cpu_req_bits_addr[0];
    end
    if (reset) begin
      wayInput <= 3'h2;
    end else if (_T_3) begin
      wayInput <= {{1'd0}, io_cpu_req_bits_way};
    end
    if (reset) begin
      replaceWayInput <= 3'h2;
    end else if (_T_3) begin
      replaceWayInput <= {{1'd0}, io_cpu_req_bits_replaceWay};
    end
    _T_54 <= decoder_io_outSignals_8;
    _T_57 <= decoder_io_outSignals_8;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_60 & _T_62) begin
          $fwrite(32'h80000002,"Replacement in Set: %d, Way: %d, Addr: %d\n",set,way,addr_reg); // @[Gem5CacheLogic.scala 461:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Gem5CacheLogic_3(
  input         clock,
  input         reset,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [27:0] io_cpu_req_bits_command,
  input  [1:0]  io_cpu_req_bits_way,
  input  [1:0]  io_cpu_req_bits_replaceWay,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_iswrite,
  output [1:0]  io_cpu_resp_bits_way,
  output        io_metaMem_write_valid,
  output [1:0]  io_metaMem_write_bits_bank,
  output        io_metaMem_write_bits_address,
  output [30:0] io_metaMem_write_bits_inputValue_0_tag,
  output [30:0] io_metaMem_write_bits_inputValue_1_tag,
  output        io_validTagBits_write_valid,
  output [63:0] io_validTagBits_write_bits_addr,
  output        io_validTagBits_write_bits_value,
  output        io_validTagBits_read_in_valid,
  output [63:0] io_validTagBits_read_in_bits_addr,
  input         io_validTagBits_read_out_0,
  input         io_validTagBits_read_out_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [27:0] decoder_io_inAction; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_7; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_8; // @[Gem5CacheLogic.scala 188:23]
  wire  emptyLine_io_data_0; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_data_1; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 359:25]
  wire [30:0] tagFinder_io_key_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_0_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_1_tag; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_0; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_1; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_value_valid; // @[Gem5CacheLogic.scala 362:25]
  wire [31:0] tagFinder_io_value_bits; // @[Gem5CacheLogic.scala 362:25]
  reg [31:0] addr_reg; // @[Gem5CacheLogic.scala 202:25]
  reg [27:0] cpu_command; // @[Gem5CacheLogic.scala 205:28]
  reg [30:0] tag; // @[Gem5CacheLogic.scala 207:20]
  reg  set; // @[Gem5CacheLogic.scala 208:20]
  reg [2:0] wayInput; // @[Gem5CacheLogic.scala 209:25]
  reg [2:0] replaceWayInput; // @[Gem5CacheLogic.scala 210:32]
  wire  _T_3 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_47 = {{1'd0}, set}; // @[Gem5CacheLogic.scala 289:41]
  wire [2:0] _T_6 = _GEN_47 * 2'h2; // @[Gem5CacheLogic.scala 289:41]
  wire  signals_2 = decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  wayInvalid = wayInput == 3'h2; // @[Gem5CacheLogic.scala 351:27]
  wire  _T_28 = ~wayInvalid; // @[Gem5CacheLogic.scala 378:14]
  wire [2:0] _GEN_15 = _T_28 ? wayInput : 3'h2; // @[Gem5CacheLogic.scala 378:26]
  wire [2:0] way = signals_2 ? replaceWayInput : _GEN_15; // @[Gem5CacheLogic.scala 376:23]
  wire [2:0] _T_8 = _T_6 + way; // @[Gem5CacheLogic.scala 289:51]
  wire  signals_1 = decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_0 = decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_23 = signals_1 & signals_0; // @[Gem5CacheLogic.scala 367:37]
  wire  _T_24 = signals_2 | _T_23; // @[Gem5CacheLogic.scala 367:21]
  wire [2:0] _GEN_14 = _T_24 ? _T_6 : 3'h0; // @[Gem5CacheLogic.scala 367:53]
  wire [7:0] _T_29 = 8'h1 << way; // @[Gem5CacheLogic.scala 338:34]
  wire  signals_4 = decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_3 = decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire [31:0] _T_47 = tagFinder_io_value_valid ? tagFinder_io_value_bits : 32'h2; // @[Gem5CacheLogic.scala 424:25]
  wire [2:0] _GEN_41 = signals_2 ? way : 3'h2; // @[Gem5CacheLogic.scala 425:28]
  wire [31:0] _GEN_43 = _T_23 ? _T_47 : {{29'd0}, _GEN_41}; // @[Gem5CacheLogic.scala 423:39]
  wire  signals_5 = decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_6 = decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_52 = ~signals_6; // @[Gem5CacheLogic.scala 446:50]
  reg  _T_54; // @[Gem5CacheLogic.scala 455:38]
  reg  _T_57; // @[Gem5CacheLogic.scala 456:81]
  wire  _T_59 = ~emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 460:26]
  wire  _T_60 = signals_2 & _T_59; // @[Gem5CacheLogic.scala 460:23]
  wire  _T_62 = ~reset; // @[Gem5CacheLogic.scala 461:13]
  wire [2:0] targetWayWire = _GEN_43[2:0]; // @[Gem5CacheLogic.scala 424:19 Gem5CacheLogic.scala 426:19]
  Decoder decoder ( // @[Gem5CacheLogic.scala 188:23]
    .io_inAction(decoder_io_inAction),
    .io_outSignals_0(decoder_io_outSignals_0),
    .io_outSignals_1(decoder_io_outSignals_1),
    .io_outSignals_2(decoder_io_outSignals_2),
    .io_outSignals_3(decoder_io_outSignals_3),
    .io_outSignals_4(decoder_io_outSignals_4),
    .io_outSignals_5(decoder_io_outSignals_5),
    .io_outSignals_6(decoder_io_outSignals_6),
    .io_outSignals_7(decoder_io_outSignals_7),
    .io_outSignals_8(decoder_io_outSignals_8)
  );
  FindEmptyLine emptyLine ( // @[Gem5CacheLogic.scala 359:25]
    .io_data_0(emptyLine_io_data_0),
    .io_data_1(emptyLine_io_data_1),
    .io_value_valid(emptyLine_io_value_valid)
  );
  Find tagFinder ( // @[Gem5CacheLogic.scala 362:25]
    .io_key_tag(tagFinder_io_key_tag),
    .io_data_0_tag(tagFinder_io_data_0_tag),
    .io_data_1_tag(tagFinder_io_data_1_tag),
    .io_valid_0(tagFinder_io_valid_0),
    .io_valid_1(tagFinder_io_valid_1),
    .io_value_valid(tagFinder_io_value_valid),
    .io_value_bits(tagFinder_io_value_bits)
  );
  assign io_cpu_req_ready = 1'h1; // @[Gem5CacheLogic.scala 302:20]
  assign io_cpu_resp_valid = _T_24 | _T_57; // @[Gem5CacheLogic.scala 456:24]
  assign io_cpu_resp_bits_iswrite = _T_54; // @[Gem5CacheLogic.scala 455:28]
  assign io_cpu_resp_bits_way = targetWayWire[1:0]; // @[Gem5CacheLogic.scala 453:24]
  assign io_metaMem_write_valid = signals_3 ? 1'h0 : signals_4; // @[Gem5CacheLogic.scala 346:26 Gem5CacheLogic.scala 330:19]
  assign io_metaMem_write_bits_bank = _T_29[1:0]; // @[Gem5CacheLogic.scala 338:27]
  assign io_metaMem_write_bits_address = set; // @[Gem5CacheLogic.scala 339:30]
  assign io_metaMem_write_bits_inputValue_0_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_metaMem_write_bits_inputValue_1_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_validTagBits_write_valid = signals_5 | signals_6; // @[Gem5CacheLogic.scala 445:31]
  assign io_validTagBits_write_bits_addr = {{61'd0}, _T_8}; // @[Gem5CacheLogic.scala 444:35]
  assign io_validTagBits_write_bits_value = signals_5 | _T_52; // @[Gem5CacheLogic.scala 446:36]
  assign io_validTagBits_read_in_valid = signals_2 | _T_23; // @[Gem5CacheLogic.scala 373:33]
  assign io_validTagBits_read_in_bits_addr = {{61'd0}, _GEN_14}; // @[Gem5CacheLogic.scala 368:39 Gem5CacheLogic.scala 370:39]
  assign decoder_io_inAction = cpu_command; // @[Gem5CacheLogic.scala 298:23]
  assign emptyLine_io_data_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 360:21]
  assign emptyLine_io_data_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 360:21]
  assign tagFinder_io_key_tag = tag; // @[Gem5CacheLogic.scala 363:20]
  assign tagFinder_io_data_0_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_data_1_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_valid_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 365:22]
  assign tagFinder_io_valid_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 365:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cpu_command = _RAND_1[27:0];
  _RAND_2 = {1{`RANDOM}};
  tag = _RAND_2[30:0];
  _RAND_3 = {1{`RANDOM}};
  set = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wayInput = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  replaceWayInput = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _T_54 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_57 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr_reg <= 32'h0;
    end else if (_T_3) begin
      addr_reg <= io_cpu_req_bits_addr;
    end
    if (reset) begin
      cpu_command <= 28'h0;
    end else if (_T_3) begin
      cpu_command <= io_cpu_req_bits_command;
    end
    if (reset) begin
      tag <= 31'h0;
    end else if (_T_3) begin
      tag <= io_cpu_req_bits_addr[31:1];
    end
    if (reset) begin
      set <= 1'h0;
    end else if (_T_3) begin
      set <= io_cpu_req_bits_addr[0];
    end
    if (reset) begin
      wayInput <= 3'h2;
    end else if (_T_3) begin
      wayInput <= {{1'd0}, io_cpu_req_bits_way};
    end
    if (reset) begin
      replaceWayInput <= 3'h2;
    end else if (_T_3) begin
      replaceWayInput <= {{1'd0}, io_cpu_req_bits_replaceWay};
    end
    _T_54 <= decoder_io_outSignals_8;
    _T_57 <= decoder_io_outSignals_8;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_60 & _T_62) begin
          $fwrite(32'h80000002,"Replacement in Set: %d, Way: %d, Addr: %d\n",set,way,addr_reg); // @[Gem5CacheLogic.scala 461:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Gem5CacheLogic_4(
  input         clock,
  input         reset,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [27:0] io_cpu_req_bits_command,
  input  [1:0]  io_cpu_req_bits_way,
  input  [1:0]  io_cpu_req_bits_replaceWay,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_iswrite,
  output [1:0]  io_cpu_resp_bits_way,
  output        io_metaMem_write_valid,
  output [1:0]  io_metaMem_write_bits_bank,
  output        io_metaMem_write_bits_address,
  output [30:0] io_metaMem_write_bits_inputValue_0_tag,
  output [30:0] io_metaMem_write_bits_inputValue_1_tag,
  output        io_validTagBits_write_valid,
  output [63:0] io_validTagBits_write_bits_addr,
  output        io_validTagBits_write_bits_value,
  output        io_validTagBits_read_in_valid,
  output [63:0] io_validTagBits_read_in_bits_addr,
  input         io_validTagBits_read_out_0,
  input         io_validTagBits_read_out_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [27:0] decoder_io_inAction; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_7; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_8; // @[Gem5CacheLogic.scala 188:23]
  wire  emptyLine_io_data_0; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_data_1; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 359:25]
  wire [30:0] tagFinder_io_key_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_0_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_1_tag; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_0; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_1; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_value_valid; // @[Gem5CacheLogic.scala 362:25]
  wire [31:0] tagFinder_io_value_bits; // @[Gem5CacheLogic.scala 362:25]
  reg [31:0] addr_reg; // @[Gem5CacheLogic.scala 202:25]
  reg [27:0] cpu_command; // @[Gem5CacheLogic.scala 205:28]
  reg [30:0] tag; // @[Gem5CacheLogic.scala 207:20]
  reg  set; // @[Gem5CacheLogic.scala 208:20]
  reg [2:0] wayInput; // @[Gem5CacheLogic.scala 209:25]
  reg [2:0] replaceWayInput; // @[Gem5CacheLogic.scala 210:32]
  wire  _T_3 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_47 = {{1'd0}, set}; // @[Gem5CacheLogic.scala 289:41]
  wire [2:0] _T_6 = _GEN_47 * 2'h2; // @[Gem5CacheLogic.scala 289:41]
  wire  signals_2 = decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  wayInvalid = wayInput == 3'h2; // @[Gem5CacheLogic.scala 351:27]
  wire  _T_28 = ~wayInvalid; // @[Gem5CacheLogic.scala 378:14]
  wire [2:0] _GEN_15 = _T_28 ? wayInput : 3'h2; // @[Gem5CacheLogic.scala 378:26]
  wire [2:0] way = signals_2 ? replaceWayInput : _GEN_15; // @[Gem5CacheLogic.scala 376:23]
  wire [2:0] _T_8 = _T_6 + way; // @[Gem5CacheLogic.scala 289:51]
  wire  signals_1 = decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_0 = decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_23 = signals_1 & signals_0; // @[Gem5CacheLogic.scala 367:37]
  wire  _T_24 = signals_2 | _T_23; // @[Gem5CacheLogic.scala 367:21]
  wire [2:0] _GEN_14 = _T_24 ? _T_6 : 3'h0; // @[Gem5CacheLogic.scala 367:53]
  wire [7:0] _T_29 = 8'h1 << way; // @[Gem5CacheLogic.scala 338:34]
  wire  signals_4 = decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_3 = decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire [31:0] _T_47 = tagFinder_io_value_valid ? tagFinder_io_value_bits : 32'h2; // @[Gem5CacheLogic.scala 424:25]
  wire [2:0] _GEN_41 = signals_2 ? way : 3'h2; // @[Gem5CacheLogic.scala 425:28]
  wire [31:0] _GEN_43 = _T_23 ? _T_47 : {{29'd0}, _GEN_41}; // @[Gem5CacheLogic.scala 423:39]
  wire  signals_5 = decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_6 = decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_52 = ~signals_6; // @[Gem5CacheLogic.scala 446:50]
  reg  _T_54; // @[Gem5CacheLogic.scala 455:38]
  reg  _T_57; // @[Gem5CacheLogic.scala 456:81]
  wire  _T_59 = ~emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 460:26]
  wire  _T_60 = signals_2 & _T_59; // @[Gem5CacheLogic.scala 460:23]
  wire  _T_62 = ~reset; // @[Gem5CacheLogic.scala 461:13]
  wire [2:0] targetWayWire = _GEN_43[2:0]; // @[Gem5CacheLogic.scala 424:19 Gem5CacheLogic.scala 426:19]
  Decoder decoder ( // @[Gem5CacheLogic.scala 188:23]
    .io_inAction(decoder_io_inAction),
    .io_outSignals_0(decoder_io_outSignals_0),
    .io_outSignals_1(decoder_io_outSignals_1),
    .io_outSignals_2(decoder_io_outSignals_2),
    .io_outSignals_3(decoder_io_outSignals_3),
    .io_outSignals_4(decoder_io_outSignals_4),
    .io_outSignals_5(decoder_io_outSignals_5),
    .io_outSignals_6(decoder_io_outSignals_6),
    .io_outSignals_7(decoder_io_outSignals_7),
    .io_outSignals_8(decoder_io_outSignals_8)
  );
  FindEmptyLine emptyLine ( // @[Gem5CacheLogic.scala 359:25]
    .io_data_0(emptyLine_io_data_0),
    .io_data_1(emptyLine_io_data_1),
    .io_value_valid(emptyLine_io_value_valid)
  );
  Find tagFinder ( // @[Gem5CacheLogic.scala 362:25]
    .io_key_tag(tagFinder_io_key_tag),
    .io_data_0_tag(tagFinder_io_data_0_tag),
    .io_data_1_tag(tagFinder_io_data_1_tag),
    .io_valid_0(tagFinder_io_valid_0),
    .io_valid_1(tagFinder_io_valid_1),
    .io_value_valid(tagFinder_io_value_valid),
    .io_value_bits(tagFinder_io_value_bits)
  );
  assign io_cpu_req_ready = 1'h1; // @[Gem5CacheLogic.scala 302:20]
  assign io_cpu_resp_valid = _T_24 | _T_57; // @[Gem5CacheLogic.scala 456:24]
  assign io_cpu_resp_bits_iswrite = _T_54; // @[Gem5CacheLogic.scala 455:28]
  assign io_cpu_resp_bits_way = targetWayWire[1:0]; // @[Gem5CacheLogic.scala 453:24]
  assign io_metaMem_write_valid = signals_3 ? 1'h0 : signals_4; // @[Gem5CacheLogic.scala 346:26 Gem5CacheLogic.scala 330:19]
  assign io_metaMem_write_bits_bank = _T_29[1:0]; // @[Gem5CacheLogic.scala 338:27]
  assign io_metaMem_write_bits_address = set; // @[Gem5CacheLogic.scala 339:30]
  assign io_metaMem_write_bits_inputValue_0_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_metaMem_write_bits_inputValue_1_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_validTagBits_write_valid = signals_5 | signals_6; // @[Gem5CacheLogic.scala 445:31]
  assign io_validTagBits_write_bits_addr = {{61'd0}, _T_8}; // @[Gem5CacheLogic.scala 444:35]
  assign io_validTagBits_write_bits_value = signals_5 | _T_52; // @[Gem5CacheLogic.scala 446:36]
  assign io_validTagBits_read_in_valid = signals_2 | _T_23; // @[Gem5CacheLogic.scala 373:33]
  assign io_validTagBits_read_in_bits_addr = {{61'd0}, _GEN_14}; // @[Gem5CacheLogic.scala 368:39 Gem5CacheLogic.scala 370:39]
  assign decoder_io_inAction = cpu_command; // @[Gem5CacheLogic.scala 298:23]
  assign emptyLine_io_data_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 360:21]
  assign emptyLine_io_data_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 360:21]
  assign tagFinder_io_key_tag = tag; // @[Gem5CacheLogic.scala 363:20]
  assign tagFinder_io_data_0_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_data_1_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_valid_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 365:22]
  assign tagFinder_io_valid_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 365:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cpu_command = _RAND_1[27:0];
  _RAND_2 = {1{`RANDOM}};
  tag = _RAND_2[30:0];
  _RAND_3 = {1{`RANDOM}};
  set = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wayInput = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  replaceWayInput = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _T_54 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_57 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr_reg <= 32'h0;
    end else if (_T_3) begin
      addr_reg <= io_cpu_req_bits_addr;
    end
    if (reset) begin
      cpu_command <= 28'h0;
    end else if (_T_3) begin
      cpu_command <= io_cpu_req_bits_command;
    end
    if (reset) begin
      tag <= 31'h0;
    end else if (_T_3) begin
      tag <= io_cpu_req_bits_addr[31:1];
    end
    if (reset) begin
      set <= 1'h0;
    end else if (_T_3) begin
      set <= io_cpu_req_bits_addr[0];
    end
    if (reset) begin
      wayInput <= 3'h2;
    end else if (_T_3) begin
      wayInput <= {{1'd0}, io_cpu_req_bits_way};
    end
    if (reset) begin
      replaceWayInput <= 3'h2;
    end else if (_T_3) begin
      replaceWayInput <= {{1'd0}, io_cpu_req_bits_replaceWay};
    end
    _T_54 <= decoder_io_outSignals_8;
    _T_57 <= decoder_io_outSignals_8;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_60 & _T_62) begin
          $fwrite(32'h80000002,"Replacement in Set: %d, Way: %d, Addr: %d\n",set,way,addr_reg); // @[Gem5CacheLogic.scala 461:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Gem5CacheLogic_5(
  input         clock,
  input         reset,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [27:0] io_cpu_req_bits_command,
  input  [1:0]  io_cpu_req_bits_way,
  input  [1:0]  io_cpu_req_bits_replaceWay,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_iswrite,
  output [1:0]  io_cpu_resp_bits_way,
  output        io_metaMem_write_valid,
  output [1:0]  io_metaMem_write_bits_bank,
  output        io_metaMem_write_bits_address,
  output [30:0] io_metaMem_write_bits_inputValue_0_tag,
  output [30:0] io_metaMem_write_bits_inputValue_1_tag,
  output        io_validTagBits_write_valid,
  output [63:0] io_validTagBits_write_bits_addr,
  output        io_validTagBits_write_bits_value,
  output        io_validTagBits_read_in_valid,
  output [63:0] io_validTagBits_read_in_bits_addr,
  input         io_validTagBits_read_out_0,
  input         io_validTagBits_read_out_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [27:0] decoder_io_inAction; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_7; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_8; // @[Gem5CacheLogic.scala 188:23]
  wire  emptyLine_io_data_0; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_data_1; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 359:25]
  wire [30:0] tagFinder_io_key_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_0_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_1_tag; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_0; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_1; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_value_valid; // @[Gem5CacheLogic.scala 362:25]
  wire [31:0] tagFinder_io_value_bits; // @[Gem5CacheLogic.scala 362:25]
  reg [31:0] addr_reg; // @[Gem5CacheLogic.scala 202:25]
  reg [27:0] cpu_command; // @[Gem5CacheLogic.scala 205:28]
  reg [30:0] tag; // @[Gem5CacheLogic.scala 207:20]
  reg  set; // @[Gem5CacheLogic.scala 208:20]
  reg [2:0] wayInput; // @[Gem5CacheLogic.scala 209:25]
  reg [2:0] replaceWayInput; // @[Gem5CacheLogic.scala 210:32]
  wire  _T_3 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_47 = {{1'd0}, set}; // @[Gem5CacheLogic.scala 289:41]
  wire [2:0] _T_6 = _GEN_47 * 2'h2; // @[Gem5CacheLogic.scala 289:41]
  wire  signals_2 = decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  wayInvalid = wayInput == 3'h2; // @[Gem5CacheLogic.scala 351:27]
  wire  _T_28 = ~wayInvalid; // @[Gem5CacheLogic.scala 378:14]
  wire [2:0] _GEN_15 = _T_28 ? wayInput : 3'h2; // @[Gem5CacheLogic.scala 378:26]
  wire [2:0] way = signals_2 ? replaceWayInput : _GEN_15; // @[Gem5CacheLogic.scala 376:23]
  wire [2:0] _T_8 = _T_6 + way; // @[Gem5CacheLogic.scala 289:51]
  wire  signals_1 = decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_0 = decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_23 = signals_1 & signals_0; // @[Gem5CacheLogic.scala 367:37]
  wire  _T_24 = signals_2 | _T_23; // @[Gem5CacheLogic.scala 367:21]
  wire [2:0] _GEN_14 = _T_24 ? _T_6 : 3'h0; // @[Gem5CacheLogic.scala 367:53]
  wire [7:0] _T_29 = 8'h1 << way; // @[Gem5CacheLogic.scala 338:34]
  wire  signals_4 = decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_3 = decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire [31:0] _T_47 = tagFinder_io_value_valid ? tagFinder_io_value_bits : 32'h2; // @[Gem5CacheLogic.scala 424:25]
  wire [2:0] _GEN_41 = signals_2 ? way : 3'h2; // @[Gem5CacheLogic.scala 425:28]
  wire [31:0] _GEN_43 = _T_23 ? _T_47 : {{29'd0}, _GEN_41}; // @[Gem5CacheLogic.scala 423:39]
  wire  signals_5 = decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_6 = decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_52 = ~signals_6; // @[Gem5CacheLogic.scala 446:50]
  reg  _T_54; // @[Gem5CacheLogic.scala 455:38]
  reg  _T_57; // @[Gem5CacheLogic.scala 456:81]
  wire  _T_59 = ~emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 460:26]
  wire  _T_60 = signals_2 & _T_59; // @[Gem5CacheLogic.scala 460:23]
  wire  _T_62 = ~reset; // @[Gem5CacheLogic.scala 461:13]
  wire [2:0] targetWayWire = _GEN_43[2:0]; // @[Gem5CacheLogic.scala 424:19 Gem5CacheLogic.scala 426:19]
  Decoder decoder ( // @[Gem5CacheLogic.scala 188:23]
    .io_inAction(decoder_io_inAction),
    .io_outSignals_0(decoder_io_outSignals_0),
    .io_outSignals_1(decoder_io_outSignals_1),
    .io_outSignals_2(decoder_io_outSignals_2),
    .io_outSignals_3(decoder_io_outSignals_3),
    .io_outSignals_4(decoder_io_outSignals_4),
    .io_outSignals_5(decoder_io_outSignals_5),
    .io_outSignals_6(decoder_io_outSignals_6),
    .io_outSignals_7(decoder_io_outSignals_7),
    .io_outSignals_8(decoder_io_outSignals_8)
  );
  FindEmptyLine emptyLine ( // @[Gem5CacheLogic.scala 359:25]
    .io_data_0(emptyLine_io_data_0),
    .io_data_1(emptyLine_io_data_1),
    .io_value_valid(emptyLine_io_value_valid)
  );
  Find tagFinder ( // @[Gem5CacheLogic.scala 362:25]
    .io_key_tag(tagFinder_io_key_tag),
    .io_data_0_tag(tagFinder_io_data_0_tag),
    .io_data_1_tag(tagFinder_io_data_1_tag),
    .io_valid_0(tagFinder_io_valid_0),
    .io_valid_1(tagFinder_io_valid_1),
    .io_value_valid(tagFinder_io_value_valid),
    .io_value_bits(tagFinder_io_value_bits)
  );
  assign io_cpu_req_ready = 1'h1; // @[Gem5CacheLogic.scala 302:20]
  assign io_cpu_resp_valid = _T_24 | _T_57; // @[Gem5CacheLogic.scala 456:24]
  assign io_cpu_resp_bits_iswrite = _T_54; // @[Gem5CacheLogic.scala 455:28]
  assign io_cpu_resp_bits_way = targetWayWire[1:0]; // @[Gem5CacheLogic.scala 453:24]
  assign io_metaMem_write_valid = signals_3 ? 1'h0 : signals_4; // @[Gem5CacheLogic.scala 346:26 Gem5CacheLogic.scala 330:19]
  assign io_metaMem_write_bits_bank = _T_29[1:0]; // @[Gem5CacheLogic.scala 338:27]
  assign io_metaMem_write_bits_address = set; // @[Gem5CacheLogic.scala 339:30]
  assign io_metaMem_write_bits_inputValue_0_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_metaMem_write_bits_inputValue_1_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_validTagBits_write_valid = signals_5 | signals_6; // @[Gem5CacheLogic.scala 445:31]
  assign io_validTagBits_write_bits_addr = {{61'd0}, _T_8}; // @[Gem5CacheLogic.scala 444:35]
  assign io_validTagBits_write_bits_value = signals_5 | _T_52; // @[Gem5CacheLogic.scala 446:36]
  assign io_validTagBits_read_in_valid = signals_2 | _T_23; // @[Gem5CacheLogic.scala 373:33]
  assign io_validTagBits_read_in_bits_addr = {{61'd0}, _GEN_14}; // @[Gem5CacheLogic.scala 368:39 Gem5CacheLogic.scala 370:39]
  assign decoder_io_inAction = cpu_command; // @[Gem5CacheLogic.scala 298:23]
  assign emptyLine_io_data_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 360:21]
  assign emptyLine_io_data_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 360:21]
  assign tagFinder_io_key_tag = tag; // @[Gem5CacheLogic.scala 363:20]
  assign tagFinder_io_data_0_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_data_1_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_valid_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 365:22]
  assign tagFinder_io_valid_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 365:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cpu_command = _RAND_1[27:0];
  _RAND_2 = {1{`RANDOM}};
  tag = _RAND_2[30:0];
  _RAND_3 = {1{`RANDOM}};
  set = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wayInput = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  replaceWayInput = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _T_54 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_57 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr_reg <= 32'h0;
    end else if (_T_3) begin
      addr_reg <= io_cpu_req_bits_addr;
    end
    if (reset) begin
      cpu_command <= 28'h0;
    end else if (_T_3) begin
      cpu_command <= io_cpu_req_bits_command;
    end
    if (reset) begin
      tag <= 31'h0;
    end else if (_T_3) begin
      tag <= io_cpu_req_bits_addr[31:1];
    end
    if (reset) begin
      set <= 1'h0;
    end else if (_T_3) begin
      set <= io_cpu_req_bits_addr[0];
    end
    if (reset) begin
      wayInput <= 3'h2;
    end else if (_T_3) begin
      wayInput <= {{1'd0}, io_cpu_req_bits_way};
    end
    if (reset) begin
      replaceWayInput <= 3'h2;
    end else if (_T_3) begin
      replaceWayInput <= {{1'd0}, io_cpu_req_bits_replaceWay};
    end
    _T_54 <= decoder_io_outSignals_8;
    _T_57 <= decoder_io_outSignals_8;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_60 & _T_62) begin
          $fwrite(32'h80000002,"Replacement in Set: %d, Way: %d, Addr: %d\n",set,way,addr_reg); // @[Gem5CacheLogic.scala 461:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Gem5CacheLogic_6(
  input         clock,
  input         reset,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [27:0] io_cpu_req_bits_command,
  input  [1:0]  io_cpu_req_bits_way,
  input  [1:0]  io_cpu_req_bits_replaceWay,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_iswrite,
  output [1:0]  io_cpu_resp_bits_way,
  output        io_metaMem_write_valid,
  output [1:0]  io_metaMem_write_bits_bank,
  output        io_metaMem_write_bits_address,
  output [30:0] io_metaMem_write_bits_inputValue_0_tag,
  output [30:0] io_metaMem_write_bits_inputValue_1_tag,
  output        io_validTagBits_write_valid,
  output [63:0] io_validTagBits_write_bits_addr,
  output        io_validTagBits_write_bits_value,
  output        io_validTagBits_read_in_valid,
  output [63:0] io_validTagBits_read_in_bits_addr,
  input         io_validTagBits_read_out_0,
  input         io_validTagBits_read_out_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [27:0] decoder_io_inAction; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_7; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_8; // @[Gem5CacheLogic.scala 188:23]
  wire  emptyLine_io_data_0; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_data_1; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 359:25]
  wire [30:0] tagFinder_io_key_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_0_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_1_tag; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_0; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_1; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_value_valid; // @[Gem5CacheLogic.scala 362:25]
  wire [31:0] tagFinder_io_value_bits; // @[Gem5CacheLogic.scala 362:25]
  reg [31:0] addr_reg; // @[Gem5CacheLogic.scala 202:25]
  reg [27:0] cpu_command; // @[Gem5CacheLogic.scala 205:28]
  reg [30:0] tag; // @[Gem5CacheLogic.scala 207:20]
  reg  set; // @[Gem5CacheLogic.scala 208:20]
  reg [2:0] wayInput; // @[Gem5CacheLogic.scala 209:25]
  reg [2:0] replaceWayInput; // @[Gem5CacheLogic.scala 210:32]
  wire  _T_3 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_47 = {{1'd0}, set}; // @[Gem5CacheLogic.scala 289:41]
  wire [2:0] _T_6 = _GEN_47 * 2'h2; // @[Gem5CacheLogic.scala 289:41]
  wire  signals_2 = decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  wayInvalid = wayInput == 3'h2; // @[Gem5CacheLogic.scala 351:27]
  wire  _T_28 = ~wayInvalid; // @[Gem5CacheLogic.scala 378:14]
  wire [2:0] _GEN_15 = _T_28 ? wayInput : 3'h2; // @[Gem5CacheLogic.scala 378:26]
  wire [2:0] way = signals_2 ? replaceWayInput : _GEN_15; // @[Gem5CacheLogic.scala 376:23]
  wire [2:0] _T_8 = _T_6 + way; // @[Gem5CacheLogic.scala 289:51]
  wire  signals_1 = decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_0 = decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_23 = signals_1 & signals_0; // @[Gem5CacheLogic.scala 367:37]
  wire  _T_24 = signals_2 | _T_23; // @[Gem5CacheLogic.scala 367:21]
  wire [2:0] _GEN_14 = _T_24 ? _T_6 : 3'h0; // @[Gem5CacheLogic.scala 367:53]
  wire [7:0] _T_29 = 8'h1 << way; // @[Gem5CacheLogic.scala 338:34]
  wire  signals_4 = decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_3 = decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire [31:0] _T_47 = tagFinder_io_value_valid ? tagFinder_io_value_bits : 32'h2; // @[Gem5CacheLogic.scala 424:25]
  wire [2:0] _GEN_41 = signals_2 ? way : 3'h2; // @[Gem5CacheLogic.scala 425:28]
  wire [31:0] _GEN_43 = _T_23 ? _T_47 : {{29'd0}, _GEN_41}; // @[Gem5CacheLogic.scala 423:39]
  wire  signals_5 = decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_6 = decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_52 = ~signals_6; // @[Gem5CacheLogic.scala 446:50]
  reg  _T_54; // @[Gem5CacheLogic.scala 455:38]
  reg  _T_57; // @[Gem5CacheLogic.scala 456:81]
  wire  _T_59 = ~emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 460:26]
  wire  _T_60 = signals_2 & _T_59; // @[Gem5CacheLogic.scala 460:23]
  wire  _T_62 = ~reset; // @[Gem5CacheLogic.scala 461:13]
  wire [2:0] targetWayWire = _GEN_43[2:0]; // @[Gem5CacheLogic.scala 424:19 Gem5CacheLogic.scala 426:19]
  Decoder decoder ( // @[Gem5CacheLogic.scala 188:23]
    .io_inAction(decoder_io_inAction),
    .io_outSignals_0(decoder_io_outSignals_0),
    .io_outSignals_1(decoder_io_outSignals_1),
    .io_outSignals_2(decoder_io_outSignals_2),
    .io_outSignals_3(decoder_io_outSignals_3),
    .io_outSignals_4(decoder_io_outSignals_4),
    .io_outSignals_5(decoder_io_outSignals_5),
    .io_outSignals_6(decoder_io_outSignals_6),
    .io_outSignals_7(decoder_io_outSignals_7),
    .io_outSignals_8(decoder_io_outSignals_8)
  );
  FindEmptyLine emptyLine ( // @[Gem5CacheLogic.scala 359:25]
    .io_data_0(emptyLine_io_data_0),
    .io_data_1(emptyLine_io_data_1),
    .io_value_valid(emptyLine_io_value_valid)
  );
  Find tagFinder ( // @[Gem5CacheLogic.scala 362:25]
    .io_key_tag(tagFinder_io_key_tag),
    .io_data_0_tag(tagFinder_io_data_0_tag),
    .io_data_1_tag(tagFinder_io_data_1_tag),
    .io_valid_0(tagFinder_io_valid_0),
    .io_valid_1(tagFinder_io_valid_1),
    .io_value_valid(tagFinder_io_value_valid),
    .io_value_bits(tagFinder_io_value_bits)
  );
  assign io_cpu_req_ready = 1'h1; // @[Gem5CacheLogic.scala 302:20]
  assign io_cpu_resp_valid = _T_24 | _T_57; // @[Gem5CacheLogic.scala 456:24]
  assign io_cpu_resp_bits_iswrite = _T_54; // @[Gem5CacheLogic.scala 455:28]
  assign io_cpu_resp_bits_way = targetWayWire[1:0]; // @[Gem5CacheLogic.scala 453:24]
  assign io_metaMem_write_valid = signals_3 ? 1'h0 : signals_4; // @[Gem5CacheLogic.scala 346:26 Gem5CacheLogic.scala 330:19]
  assign io_metaMem_write_bits_bank = _T_29[1:0]; // @[Gem5CacheLogic.scala 338:27]
  assign io_metaMem_write_bits_address = set; // @[Gem5CacheLogic.scala 339:30]
  assign io_metaMem_write_bits_inputValue_0_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_metaMem_write_bits_inputValue_1_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_validTagBits_write_valid = signals_5 | signals_6; // @[Gem5CacheLogic.scala 445:31]
  assign io_validTagBits_write_bits_addr = {{61'd0}, _T_8}; // @[Gem5CacheLogic.scala 444:35]
  assign io_validTagBits_write_bits_value = signals_5 | _T_52; // @[Gem5CacheLogic.scala 446:36]
  assign io_validTagBits_read_in_valid = signals_2 | _T_23; // @[Gem5CacheLogic.scala 373:33]
  assign io_validTagBits_read_in_bits_addr = {{61'd0}, _GEN_14}; // @[Gem5CacheLogic.scala 368:39 Gem5CacheLogic.scala 370:39]
  assign decoder_io_inAction = cpu_command; // @[Gem5CacheLogic.scala 298:23]
  assign emptyLine_io_data_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 360:21]
  assign emptyLine_io_data_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 360:21]
  assign tagFinder_io_key_tag = tag; // @[Gem5CacheLogic.scala 363:20]
  assign tagFinder_io_data_0_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_data_1_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_valid_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 365:22]
  assign tagFinder_io_valid_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 365:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cpu_command = _RAND_1[27:0];
  _RAND_2 = {1{`RANDOM}};
  tag = _RAND_2[30:0];
  _RAND_3 = {1{`RANDOM}};
  set = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wayInput = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  replaceWayInput = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _T_54 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_57 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr_reg <= 32'h0;
    end else if (_T_3) begin
      addr_reg <= io_cpu_req_bits_addr;
    end
    if (reset) begin
      cpu_command <= 28'h0;
    end else if (_T_3) begin
      cpu_command <= io_cpu_req_bits_command;
    end
    if (reset) begin
      tag <= 31'h0;
    end else if (_T_3) begin
      tag <= io_cpu_req_bits_addr[31:1];
    end
    if (reset) begin
      set <= 1'h0;
    end else if (_T_3) begin
      set <= io_cpu_req_bits_addr[0];
    end
    if (reset) begin
      wayInput <= 3'h2;
    end else if (_T_3) begin
      wayInput <= {{1'd0}, io_cpu_req_bits_way};
    end
    if (reset) begin
      replaceWayInput <= 3'h2;
    end else if (_T_3) begin
      replaceWayInput <= {{1'd0}, io_cpu_req_bits_replaceWay};
    end
    _T_54 <= decoder_io_outSignals_8;
    _T_57 <= decoder_io_outSignals_8;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_60 & _T_62) begin
          $fwrite(32'h80000002,"Replacement in Set: %d, Way: %d, Addr: %d\n",set,way,addr_reg); // @[Gem5CacheLogic.scala 461:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Gem5CacheLogic_7(
  input         clock,
  input         reset,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [63:0] io_cpu_req_bits_data,
  input  [27:0] io_cpu_req_bits_command,
  input  [1:0]  io_cpu_req_bits_way,
  input  [1:0]  io_cpu_req_bits_replaceWay,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_iswrite,
  output [1:0]  io_cpu_resp_bits_way,
  output        io_metaMem_write_valid,
  output [1:0]  io_metaMem_write_bits_bank,
  output        io_metaMem_write_bits_address,
  output [30:0] io_metaMem_write_bits_inputValue_0_tag,
  output [30:0] io_metaMem_write_bits_inputValue_1_tag,
  output        io_dataMem_write_valid,
  output [31:0] io_dataMem_write_bits_address,
  output [63:0] io_dataMem_write_bits_inputValue_0,
  output        io_validTagBits_write_valid,
  output [63:0] io_validTagBits_write_bits_addr,
  output        io_validTagBits_write_bits_value,
  output        io_validTagBits_read_in_valid,
  output [63:0] io_validTagBits_read_in_bits_addr,
  input         io_validTagBits_read_out_0,
  input         io_validTagBits_read_out_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire [27:0] decoder_io_inAction; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_7; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_8; // @[Gem5CacheLogic.scala 188:23]
  wire  emptyLine_io_data_0; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_data_1; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 359:25]
  wire [30:0] tagFinder_io_key_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_0_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [30:0] tagFinder_io_data_1_tag; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_0; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_1; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_value_valid; // @[Gem5CacheLogic.scala 362:25]
  wire [31:0] tagFinder_io_value_bits; // @[Gem5CacheLogic.scala 362:25]
  reg [31:0] addr_reg; // @[Gem5CacheLogic.scala 202:25]
  reg [63:0] cpu_data; // @[Gem5CacheLogic.scala 203:25]
  reg [27:0] cpu_command; // @[Gem5CacheLogic.scala 205:28]
  reg [30:0] tag; // @[Gem5CacheLogic.scala 207:20]
  reg  set; // @[Gem5CacheLogic.scala 208:20]
  reg [2:0] wayInput; // @[Gem5CacheLogic.scala 209:25]
  reg [2:0] replaceWayInput; // @[Gem5CacheLogic.scala 210:32]
  wire  _T_3 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_47 = {{1'd0}, set}; // @[Gem5CacheLogic.scala 289:41]
  wire [2:0] _T_6 = _GEN_47 * 2'h2; // @[Gem5CacheLogic.scala 289:41]
  wire  signals_2 = decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  wayInvalid = wayInput == 3'h2; // @[Gem5CacheLogic.scala 351:27]
  wire  _T_28 = ~wayInvalid; // @[Gem5CacheLogic.scala 378:14]
  wire [2:0] _GEN_15 = _T_28 ? wayInput : 3'h2; // @[Gem5CacheLogic.scala 378:26]
  wire [2:0] way = signals_2 ? replaceWayInput : _GEN_15; // @[Gem5CacheLogic.scala 376:23]
  wire [2:0] _T_8 = _T_6 + way; // @[Gem5CacheLogic.scala 289:51]
  wire  signals_1 = decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_0 = decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_23 = signals_1 & signals_0; // @[Gem5CacheLogic.scala 367:37]
  wire  _T_24 = signals_2 | _T_23; // @[Gem5CacheLogic.scala 367:21]
  wire [2:0] _GEN_14 = _T_24 ? _T_6 : 3'h0; // @[Gem5CacheLogic.scala 367:53]
  wire [7:0] _T_29 = 8'h1 << way; // @[Gem5CacheLogic.scala 338:34]
  wire  signals_4 = decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_3 = decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire [31:0] _T_47 = tagFinder_io_value_valid ? tagFinder_io_value_bits : 32'h2; // @[Gem5CacheLogic.scala 424:25]
  wire [2:0] _GEN_41 = signals_2 ? way : 3'h2; // @[Gem5CacheLogic.scala 425:28]
  wire [31:0] _GEN_43 = _T_23 ? _T_47 : {{29'd0}, _GEN_41}; // @[Gem5CacheLogic.scala 423:39]
  wire  signals_5 = decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_6 = decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_52 = ~signals_6; // @[Gem5CacheLogic.scala 446:50]
  reg  _T_54; // @[Gem5CacheLogic.scala 455:38]
  reg  _T_57; // @[Gem5CacheLogic.scala 456:81]
  wire  _T_59 = ~emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 460:26]
  wire  _T_60 = signals_2 & _T_59; // @[Gem5CacheLogic.scala 460:23]
  wire  _T_62 = ~reset; // @[Gem5CacheLogic.scala 461:13]
  wire [2:0] targetWayWire = _GEN_43[2:0]; // @[Gem5CacheLogic.scala 424:19 Gem5CacheLogic.scala 426:19]
  Decoder decoder ( // @[Gem5CacheLogic.scala 188:23]
    .io_inAction(decoder_io_inAction),
    .io_outSignals_0(decoder_io_outSignals_0),
    .io_outSignals_1(decoder_io_outSignals_1),
    .io_outSignals_2(decoder_io_outSignals_2),
    .io_outSignals_3(decoder_io_outSignals_3),
    .io_outSignals_4(decoder_io_outSignals_4),
    .io_outSignals_5(decoder_io_outSignals_5),
    .io_outSignals_6(decoder_io_outSignals_6),
    .io_outSignals_7(decoder_io_outSignals_7),
    .io_outSignals_8(decoder_io_outSignals_8)
  );
  FindEmptyLine emptyLine ( // @[Gem5CacheLogic.scala 359:25]
    .io_data_0(emptyLine_io_data_0),
    .io_data_1(emptyLine_io_data_1),
    .io_value_valid(emptyLine_io_value_valid)
  );
  Find tagFinder ( // @[Gem5CacheLogic.scala 362:25]
    .io_key_tag(tagFinder_io_key_tag),
    .io_data_0_tag(tagFinder_io_data_0_tag),
    .io_data_1_tag(tagFinder_io_data_1_tag),
    .io_valid_0(tagFinder_io_valid_0),
    .io_valid_1(tagFinder_io_valid_1),
    .io_value_valid(tagFinder_io_value_valid),
    .io_value_bits(tagFinder_io_value_bits)
  );
  assign io_cpu_req_ready = 1'h1; // @[Gem5CacheLogic.scala 302:20]
  assign io_cpu_resp_valid = _T_24 | _T_57; // @[Gem5CacheLogic.scala 456:24]
  assign io_cpu_resp_bits_iswrite = _T_54; // @[Gem5CacheLogic.scala 455:28]
  assign io_cpu_resp_bits_way = targetWayWire[1:0]; // @[Gem5CacheLogic.scala 453:24]
  assign io_metaMem_write_valid = signals_3 ? 1'h0 : signals_4; // @[Gem5CacheLogic.scala 346:26 Gem5CacheLogic.scala 330:19]
  assign io_metaMem_write_bits_bank = _T_29[1:0]; // @[Gem5CacheLogic.scala 338:27]
  assign io_metaMem_write_bits_address = set; // @[Gem5CacheLogic.scala 339:30]
  assign io_metaMem_write_bits_inputValue_0_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_metaMem_write_bits_inputValue_1_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_dataMem_write_valid = decoder_io_outSignals_7; // @[Gem5CacheLogic.scala 347:26 Gem5CacheLogic.scala 330:19]
  assign io_dataMem_write_bits_address = {{29'd0}, _T_8}; // @[Gem5CacheLogic.scala 334:30]
  assign io_dataMem_write_bits_inputValue_0 = cpu_data; // @[Gem5CacheLogic.scala 397:38]
  assign io_validTagBits_write_valid = signals_5 | signals_6; // @[Gem5CacheLogic.scala 445:31]
  assign io_validTagBits_write_bits_addr = {{61'd0}, _T_8}; // @[Gem5CacheLogic.scala 444:35]
  assign io_validTagBits_write_bits_value = signals_5 | _T_52; // @[Gem5CacheLogic.scala 446:36]
  assign io_validTagBits_read_in_valid = signals_2 | _T_23; // @[Gem5CacheLogic.scala 373:33]
  assign io_validTagBits_read_in_bits_addr = {{61'd0}, _GEN_14}; // @[Gem5CacheLogic.scala 368:39 Gem5CacheLogic.scala 370:39]
  assign decoder_io_inAction = cpu_command; // @[Gem5CacheLogic.scala 298:23]
  assign emptyLine_io_data_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 360:21]
  assign emptyLine_io_data_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 360:21]
  assign tagFinder_io_key_tag = tag; // @[Gem5CacheLogic.scala 363:20]
  assign tagFinder_io_data_0_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_data_1_tag = 31'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_valid_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 365:22]
  assign tagFinder_io_valid_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 365:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  cpu_data = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  cpu_command = _RAND_2[27:0];
  _RAND_3 = {1{`RANDOM}};
  tag = _RAND_3[30:0];
  _RAND_4 = {1{`RANDOM}};
  set = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wayInput = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  replaceWayInput = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _T_54 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_57 = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr_reg <= 32'h0;
    end else if (_T_3) begin
      addr_reg <= io_cpu_req_bits_addr;
    end
    if (reset) begin
      cpu_data <= 64'h0;
    end else if (_T_3) begin
      cpu_data <= io_cpu_req_bits_data;
    end
    if (reset) begin
      cpu_command <= 28'h0;
    end else if (_T_3) begin
      cpu_command <= io_cpu_req_bits_command;
    end
    if (reset) begin
      tag <= 31'h0;
    end else if (_T_3) begin
      tag <= io_cpu_req_bits_addr[31:1];
    end
    if (reset) begin
      set <= 1'h0;
    end else if (_T_3) begin
      set <= io_cpu_req_bits_addr[0];
    end
    if (reset) begin
      wayInput <= 3'h2;
    end else if (_T_3) begin
      wayInput <= {{1'd0}, io_cpu_req_bits_way};
    end
    if (reset) begin
      replaceWayInput <= 3'h2;
    end else if (_T_3) begin
      replaceWayInput <= {{1'd0}, io_cpu_req_bits_replaceWay};
    end
    _T_54 <= decoder_io_outSignals_8;
    _T_57 <= decoder_io_outSignals_8;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_60 & _T_62) begin
          $fwrite(32'h80000002,"Replacement in Set: %d, Way: %d, Addr: %d\n",set,way,addr_reg); // @[Gem5CacheLogic.scala 461:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module FindMultiLine(
  input  [30:0] io_key_tag,
  input  [30:0] io_data_0_tag,
  input  [30:0] io_data_1_tag,
  output        io_value_bits_0,
  output        io_value_bits_1
);
  wire  _T = io_data_0_tag == io_key_tag; // @[elements.scala 54:54]
  wire  _T_1 = io_data_1_tag == io_key_tag; // @[elements.scala 54:54]
  wire [1:0] bitmap = {_T_1,_T}; // @[Cat.scala 29:58]
  assign io_value_bits_0 = bitmap[0]; // @[elements.scala 57:19]
  assign io_value_bits_1 = bitmap[1]; // @[elements.scala 57:19]
endmodule
module ProbeUnit(
  input         clock,
  input         reset,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [27:0] io_cpu_req_bits_command,
  output        io_cpu_resp_valid,
  output [1:0]  io_cpu_resp_bits_way,
  output        io_cpu_multiWay_valid,
  output [1:0]  io_cpu_multiWay_bits_way_0,
  output [1:0]  io_cpu_multiWay_bits_way_1,
  output [31:0] io_cpu_multiWay_bits_addr,
  output        io_metaMem_read_in_valid,
  output        io_metaMem_read_in_bits_address,
  input  [30:0] io_metaMem_read_outputValue_0_tag,
  input  [30:0] io_metaMem_read_outputValue_1_tag,
  output        io_validTagBits_write_valid,
  output [63:0] io_validTagBits_write_bits_addr,
  output        io_validTagBits_write_bits_value,
  output        io_validTagBits_read_in_valid,
  output [63:0] io_validTagBits_read_in_bits_addr,
  input         io_validTagBits_read_out_0,
  input         io_validTagBits_read_out_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [27:0] decoder_io_inAction; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_0; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_1; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_2; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_3; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_4; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_5; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_6; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_7; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_8; // @[ProbeUnit.scala 48:23]
  wire  emptyLine_io_data_0; // @[ProbeUnit.scala 217:25]
  wire  emptyLine_io_data_1; // @[ProbeUnit.scala 217:25]
  wire  emptyLine_io_value_valid; // @[ProbeUnit.scala 217:25]
  wire [30:0] multiTagFinder_io_key_tag; // @[ProbeUnit.scala 220:30]
  wire [30:0] multiTagFinder_io_data_0_tag; // @[ProbeUnit.scala 220:30]
  wire [30:0] multiTagFinder_io_data_1_tag; // @[ProbeUnit.scala 220:30]
  wire  multiTagFinder_io_value_bits_0; // @[ProbeUnit.scala 220:30]
  wire  multiTagFinder_io_value_bits_1; // @[ProbeUnit.scala 220:30]
  wire [30:0] tagFinder_io_key_tag; // @[ProbeUnit.scala 221:25]
  wire [30:0] tagFinder_io_data_0_tag; // @[ProbeUnit.scala 221:25]
  wire [30:0] tagFinder_io_data_1_tag; // @[ProbeUnit.scala 221:25]
  wire  tagFinder_io_valid_0; // @[ProbeUnit.scala 221:25]
  wire  tagFinder_io_valid_1; // @[ProbeUnit.scala 221:25]
  wire  tagFinder_io_value_valid; // @[ProbeUnit.scala 221:25]
  wire [31:0] tagFinder_io_value_bits; // @[ProbeUnit.scala 221:25]
  reg [31:0] addr_reg; // @[ProbeUnit.scala 61:25]
  reg [27:0] cpu_command; // @[ProbeUnit.scala 64:28]
  reg [30:0] tag; // @[ProbeUnit.scala 66:20]
  reg  set; // @[ProbeUnit.scala 67:20]
  reg [2:0] wayInput; // @[ProbeUnit.scala 68:25]
  reg [2:0] replaceWayInput; // @[ProbeUnit.scala 69:32]
  wire  _T_4 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_47 = {{1'd0}, set}; // @[ProbeUnit.scala 146:41]
  wire [2:0] _T_8 = _GEN_47 * 2'h2; // @[ProbeUnit.scala 146:41]
  wire  signals_2 = decoder_io_outSignals_2; // @[ProbeUnit.scala 87:21 ProbeUnit.scala 156:11]
  wire  wayInvalid = wayInput == 3'h2; // @[ProbeUnit.scala 209:27]
  wire  _T_30 = ~wayInvalid; // @[ProbeUnit.scala 245:14]
  wire [2:0] _GEN_15 = _T_30 ? wayInput : 3'h2; // @[ProbeUnit.scala 245:26]
  wire [2:0] way = signals_2 ? replaceWayInput : _GEN_15; // @[ProbeUnit.scala 243:23]
  wire [2:0] _T_10 = _T_8 + way; // @[ProbeUnit.scala 146:51]
  wire  signals_1 = decoder_io_outSignals_1; // @[ProbeUnit.scala 87:21 ProbeUnit.scala 156:11]
  wire  signals_0 = decoder_io_outSignals_0; // @[ProbeUnit.scala 87:21 ProbeUnit.scala 156:11]
  wire  _T_25 = signals_1 & signals_0; // @[ProbeUnit.scala 234:37]
  wire  _T_26 = signals_2 | _T_25; // @[ProbeUnit.scala 234:21]
  wire [2:0] _GEN_14 = _T_26 ? _T_8 : 3'h0; // @[ProbeUnit.scala 234:53]
  wire [31:0] _T_49 = tagFinder_io_value_valid ? tagFinder_io_value_bits : 32'h2; // @[ProbeUnit.scala 287:25]
  wire [2:0] _GEN_41 = signals_2 ? way : 3'h2; // @[ProbeUnit.scala 288:28]
  wire [31:0] _GEN_42 = _T_25 ? _T_49 : {{29'd0}, _GEN_41}; // @[ProbeUnit.scala 286:39]
  wire  _T_51 = multiTagFinder_io_value_bits_0; // @[ProbeUnit.scala 294:74]
  wire [1:0] _T_52 = _T_51 ? 2'h0 : 2'h2; // @[ProbeUnit.scala 294:35]
  wire  _T_53 = multiTagFinder_io_value_bits_1; // @[ProbeUnit.scala 294:74]
  wire [1:0] _T_54 = _T_53 ? 2'h1 : 2'h2; // @[ProbeUnit.scala 294:35]
  wire  signals_5 = decoder_io_outSignals_5; // @[ProbeUnit.scala 87:21 ProbeUnit.scala 156:11]
  wire  signals_6 = decoder_io_outSignals_6; // @[ProbeUnit.scala 87:21 ProbeUnit.scala 156:11]
  wire  _T_59 = ~signals_6; // @[ProbeUnit.scala 311:50]
  wire [2:0] targetWayWire = _GEN_42[2:0]; // @[ProbeUnit.scala 287:19 ProbeUnit.scala 289:19]
  Decoder decoder ( // @[ProbeUnit.scala 48:23]
    .io_inAction(decoder_io_inAction),
    .io_outSignals_0(decoder_io_outSignals_0),
    .io_outSignals_1(decoder_io_outSignals_1),
    .io_outSignals_2(decoder_io_outSignals_2),
    .io_outSignals_3(decoder_io_outSignals_3),
    .io_outSignals_4(decoder_io_outSignals_4),
    .io_outSignals_5(decoder_io_outSignals_5),
    .io_outSignals_6(decoder_io_outSignals_6),
    .io_outSignals_7(decoder_io_outSignals_7),
    .io_outSignals_8(decoder_io_outSignals_8)
  );
  FindEmptyLine emptyLine ( // @[ProbeUnit.scala 217:25]
    .io_data_0(emptyLine_io_data_0),
    .io_data_1(emptyLine_io_data_1),
    .io_value_valid(emptyLine_io_value_valid)
  );
  FindMultiLine multiTagFinder ( // @[ProbeUnit.scala 220:30]
    .io_key_tag(multiTagFinder_io_key_tag),
    .io_data_0_tag(multiTagFinder_io_data_0_tag),
    .io_data_1_tag(multiTagFinder_io_data_1_tag),
    .io_value_bits_0(multiTagFinder_io_value_bits_0),
    .io_value_bits_1(multiTagFinder_io_value_bits_1)
  );
  Find tagFinder ( // @[ProbeUnit.scala 221:25]
    .io_key_tag(tagFinder_io_key_tag),
    .io_data_0_tag(tagFinder_io_data_0_tag),
    .io_data_1_tag(tagFinder_io_data_1_tag),
    .io_valid_0(tagFinder_io_valid_0),
    .io_valid_1(tagFinder_io_valid_1),
    .io_value_valid(tagFinder_io_value_valid),
    .io_value_bits(tagFinder_io_value_bits)
  );
  assign io_cpu_req_ready = 1'h1; // @[ProbeUnit.scala 159:20]
  assign io_cpu_resp_valid = signals_1 & signals_0; // @[ProbeUnit.scala 321:24]
  assign io_cpu_resp_bits_way = targetWayWire[1:0]; // @[ProbeUnit.scala 318:24]
  assign io_cpu_multiWay_valid = io_cpu_resp_valid; // @[ProbeUnit.scala 322:25]
  assign io_cpu_multiWay_bits_way_0 = _T_25 ? _T_52 : 2'h0; // @[ProbeUnit.scala 315:28]
  assign io_cpu_multiWay_bits_way_1 = _T_25 ? _T_54 : 2'h0; // @[ProbeUnit.scala 315:28]
  assign io_cpu_multiWay_bits_addr = addr_reg; // @[ProbeUnit.scala 316:29]
  assign io_metaMem_read_in_valid = decoder_io_outSignals_3; // @[ProbeUnit.scala 206:28 ProbeUnit.scala 172:21]
  assign io_metaMem_read_in_bits_address = set; // @[ProbeUnit.scala 181:32]
  assign io_validTagBits_write_valid = signals_5 | signals_6; // @[ProbeUnit.scala 310:31]
  assign io_validTagBits_write_bits_addr = {{61'd0}, _T_10}; // @[ProbeUnit.scala 309:35]
  assign io_validTagBits_write_bits_value = signals_5 | _T_59; // @[ProbeUnit.scala 311:36]
  assign io_validTagBits_read_in_valid = signals_2 | _T_25; // @[ProbeUnit.scala 240:33]
  assign io_validTagBits_read_in_bits_addr = {{61'd0}, _GEN_14}; // @[ProbeUnit.scala 235:39 ProbeUnit.scala 237:39]
  assign decoder_io_inAction = cpu_command; // @[ProbeUnit.scala 155:23]
  assign emptyLine_io_data_0 = io_validTagBits_read_out_0; // @[ProbeUnit.scala 218:21]
  assign emptyLine_io_data_1 = io_validTagBits_read_out_1; // @[ProbeUnit.scala 218:21]
  assign multiTagFinder_io_key_tag = tag; // @[ProbeUnit.scala 227:25]
  assign multiTagFinder_io_data_0_tag = io_metaMem_read_outputValue_0_tag; // @[ProbeUnit.scala 228:26]
  assign multiTagFinder_io_data_1_tag = io_metaMem_read_outputValue_1_tag; // @[ProbeUnit.scala 228:26]
  assign tagFinder_io_key_tag = tag; // @[ProbeUnit.scala 223:20]
  assign tagFinder_io_data_0_tag = io_metaMem_read_outputValue_0_tag; // @[ProbeUnit.scala 224:21]
  assign tagFinder_io_data_1_tag = io_metaMem_read_outputValue_1_tag; // @[ProbeUnit.scala 224:21]
  assign tagFinder_io_valid_0 = io_validTagBits_read_out_0; // @[ProbeUnit.scala 225:22]
  assign tagFinder_io_valid_1 = io_validTagBits_read_out_1; // @[ProbeUnit.scala 225:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cpu_command = _RAND_1[27:0];
  _RAND_2 = {1{`RANDOM}};
  tag = _RAND_2[30:0];
  _RAND_3 = {1{`RANDOM}};
  set = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wayInput = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  replaceWayInput = _RAND_5[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr_reg <= 32'h0;
    end else if (_T_4) begin
      addr_reg <= io_cpu_req_bits_addr;
    end
    if (reset) begin
      cpu_command <= 28'h0;
    end else if (_T_4) begin
      cpu_command <= io_cpu_req_bits_command;
    end else begin
      cpu_command <= 28'h0;
    end
    if (reset) begin
      tag <= 31'h0;
    end else if (_T_4) begin
      tag <= io_cpu_req_bits_addr[31:1];
    end
    if (reset) begin
      set <= 1'h0;
    end else if (_T_4) begin
      set <= io_cpu_req_bits_addr[0];
    end
    if (reset) begin
      wayInput <= 3'h2;
    end else if (_T_4) begin
      wayInput <= 3'h0;
    end
    if (reset) begin
      replaceWayInput <= 3'h2;
    end else if (_T_4) begin
      replaceWayInput <= 3'h0;
    end
  end
endmodule
module paralReg_1(
  input         clock,
  input         reset,
  input         io_port_0_write_valid,
  input  [63:0] io_port_0_write_bits_addr,
  input         io_port_0_write_bits_value,
  input         io_port_0_read_in_valid,
  input  [63:0] io_port_0_read_in_bits_addr,
  output        io_port_0_read_out_0,
  output        io_port_0_read_out_1,
  input         io_port_1_write_valid,
  input  [63:0] io_port_1_write_bits_addr,
  input         io_port_1_write_bits_value,
  input         io_port_1_read_in_valid,
  input  [63:0] io_port_1_read_in_bits_addr,
  output        io_port_1_read_out_0,
  output        io_port_1_read_out_1,
  input         io_port_2_write_valid,
  input  [63:0] io_port_2_write_bits_addr,
  input         io_port_2_write_bits_value,
  input         io_port_2_read_in_valid,
  input  [63:0] io_port_2_read_in_bits_addr,
  output        io_port_2_read_out_0,
  output        io_port_2_read_out_1,
  input         io_port_3_write_valid,
  input  [63:0] io_port_3_write_bits_addr,
  input         io_port_3_write_bits_value,
  input         io_port_3_read_in_valid,
  input  [63:0] io_port_3_read_in_bits_addr,
  output        io_port_3_read_out_0,
  output        io_port_3_read_out_1,
  input         io_port_4_write_valid,
  input  [63:0] io_port_4_write_bits_addr,
  input         io_port_4_write_bits_value,
  input         io_port_4_read_in_valid,
  input  [63:0] io_port_4_read_in_bits_addr,
  output        io_port_4_read_out_0,
  output        io_port_4_read_out_1,
  input         io_port_5_write_valid,
  input  [63:0] io_port_5_write_bits_addr,
  input         io_port_5_write_bits_value,
  input         io_port_5_read_in_valid,
  input  [63:0] io_port_5_read_in_bits_addr,
  output        io_port_5_read_out_0,
  output        io_port_5_read_out_1,
  input         io_port_6_write_valid,
  input  [63:0] io_port_6_write_bits_addr,
  input         io_port_6_write_bits_value,
  input         io_port_6_read_in_valid,
  input  [63:0] io_port_6_read_in_bits_addr,
  output        io_port_6_read_out_0,
  output        io_port_6_read_out_1,
  input         io_port_7_write_valid,
  input  [63:0] io_port_7_write_bits_addr,
  input         io_port_7_write_bits_value,
  input         io_port_7_read_in_valid,
  input  [63:0] io_port_7_read_in_bits_addr,
  output        io_port_7_read_out_0,
  output        io_port_7_read_out_1,
  input         io_port_8_write_valid,
  input  [63:0] io_port_8_write_bits_addr,
  input         io_port_8_write_bits_value,
  input         io_port_8_read_in_valid,
  input  [63:0] io_port_8_read_in_bits_addr,
  output        io_port_8_read_out_0,
  output        io_port_8_read_out_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  content_0; // @[elements.scala 107:26]
  reg  content_1; // @[elements.scala 107:26]
  reg  content_2; // @[elements.scala 107:26]
  reg  content_3; // @[elements.scala 107:26]
  wire [64:0] _T_1 = {{1'd0}, io_port_0_read_in_bits_addr}; // @[elements.scala 118:104]
  wire [63:0] _T_5 = io_port_0_read_in_bits_addr + 64'h1; // @[elements.scala 118:104]
  wire  _GEN_1 = 2'h1 == _T_5[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_2 = 2'h2 == _T_5[1:0] ? content_2 : _GEN_1; // @[Cat.scala 29:58]
  wire  _GEN_3 = 2'h3 == _T_5[1:0] ? content_3 : _GEN_2; // @[Cat.scala 29:58]
  wire  _GEN_5 = 2'h1 == _T_1[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_6 = 2'h2 == _T_1[1:0] ? content_2 : _GEN_5; // @[Cat.scala 29:58]
  wire  _GEN_7 = 2'h3 == _T_1[1:0] ? content_3 : _GEN_6; // @[Cat.scala 29:58]
  wire [1:0] _T_7 = {_GEN_3,_GEN_7}; // @[Cat.scala 29:58]
  wire  _GEN_10 = 2'h0 == io_port_0_write_bits_addr[1:0] ? io_port_0_write_bits_value : content_0; // @[elements.scala 124:49]
  wire  _GEN_11 = 2'h1 == io_port_0_write_bits_addr[1:0] ? io_port_0_write_bits_value : content_1; // @[elements.scala 124:49]
  wire  _GEN_12 = 2'h2 == io_port_0_write_bits_addr[1:0] ? io_port_0_write_bits_value : content_2; // @[elements.scala 124:49]
  wire  _GEN_13 = 2'h3 == io_port_0_write_bits_addr[1:0] ? io_port_0_write_bits_value : content_3; // @[elements.scala 124:49]
  wire  _GEN_14 = io_port_0_write_valid ? _GEN_10 : content_0; // @[elements.scala 123:26]
  wire  _GEN_15 = io_port_0_write_valid ? _GEN_11 : content_1; // @[elements.scala 123:26]
  wire  _GEN_16 = io_port_0_write_valid ? _GEN_12 : content_2; // @[elements.scala 123:26]
  wire  _GEN_17 = io_port_0_write_valid ? _GEN_13 : content_3; // @[elements.scala 123:26]
  wire [64:0] _T_18 = {{1'd0}, io_port_1_read_in_bits_addr}; // @[elements.scala 118:104]
  wire [63:0] _T_22 = io_port_1_read_in_bits_addr + 64'h1; // @[elements.scala 118:104]
  wire  _GEN_19 = 2'h1 == _T_22[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_20 = 2'h2 == _T_22[1:0] ? content_2 : _GEN_19; // @[Cat.scala 29:58]
  wire  _GEN_21 = 2'h3 == _T_22[1:0] ? content_3 : _GEN_20; // @[Cat.scala 29:58]
  wire  _GEN_23 = 2'h1 == _T_18[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_24 = 2'h2 == _T_18[1:0] ? content_2 : _GEN_23; // @[Cat.scala 29:58]
  wire  _GEN_25 = 2'h3 == _T_18[1:0] ? content_3 : _GEN_24; // @[Cat.scala 29:58]
  wire [1:0] _T_24 = {_GEN_21,_GEN_25}; // @[Cat.scala 29:58]
  wire  _GEN_28 = 2'h0 == io_port_1_write_bits_addr[1:0] ? io_port_1_write_bits_value : _GEN_14; // @[elements.scala 124:49]
  wire  _GEN_29 = 2'h1 == io_port_1_write_bits_addr[1:0] ? io_port_1_write_bits_value : _GEN_15; // @[elements.scala 124:49]
  wire  _GEN_30 = 2'h2 == io_port_1_write_bits_addr[1:0] ? io_port_1_write_bits_value : _GEN_16; // @[elements.scala 124:49]
  wire  _GEN_31 = 2'h3 == io_port_1_write_bits_addr[1:0] ? io_port_1_write_bits_value : _GEN_17; // @[elements.scala 124:49]
  wire  _GEN_32 = io_port_1_write_valid ? _GEN_28 : _GEN_14; // @[elements.scala 123:26]
  wire  _GEN_33 = io_port_1_write_valid ? _GEN_29 : _GEN_15; // @[elements.scala 123:26]
  wire  _GEN_34 = io_port_1_write_valid ? _GEN_30 : _GEN_16; // @[elements.scala 123:26]
  wire  _GEN_35 = io_port_1_write_valid ? _GEN_31 : _GEN_17; // @[elements.scala 123:26]
  wire [64:0] _T_35 = {{1'd0}, io_port_2_read_in_bits_addr}; // @[elements.scala 118:104]
  wire [63:0] _T_39 = io_port_2_read_in_bits_addr + 64'h1; // @[elements.scala 118:104]
  wire  _GEN_37 = 2'h1 == _T_39[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_38 = 2'h2 == _T_39[1:0] ? content_2 : _GEN_37; // @[Cat.scala 29:58]
  wire  _GEN_39 = 2'h3 == _T_39[1:0] ? content_3 : _GEN_38; // @[Cat.scala 29:58]
  wire  _GEN_41 = 2'h1 == _T_35[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_42 = 2'h2 == _T_35[1:0] ? content_2 : _GEN_41; // @[Cat.scala 29:58]
  wire  _GEN_43 = 2'h3 == _T_35[1:0] ? content_3 : _GEN_42; // @[Cat.scala 29:58]
  wire [1:0] _T_41 = {_GEN_39,_GEN_43}; // @[Cat.scala 29:58]
  wire  _GEN_46 = 2'h0 == io_port_2_write_bits_addr[1:0] ? io_port_2_write_bits_value : _GEN_32; // @[elements.scala 124:49]
  wire  _GEN_47 = 2'h1 == io_port_2_write_bits_addr[1:0] ? io_port_2_write_bits_value : _GEN_33; // @[elements.scala 124:49]
  wire  _GEN_48 = 2'h2 == io_port_2_write_bits_addr[1:0] ? io_port_2_write_bits_value : _GEN_34; // @[elements.scala 124:49]
  wire  _GEN_49 = 2'h3 == io_port_2_write_bits_addr[1:0] ? io_port_2_write_bits_value : _GEN_35; // @[elements.scala 124:49]
  wire  _GEN_50 = io_port_2_write_valid ? _GEN_46 : _GEN_32; // @[elements.scala 123:26]
  wire  _GEN_51 = io_port_2_write_valid ? _GEN_47 : _GEN_33; // @[elements.scala 123:26]
  wire  _GEN_52 = io_port_2_write_valid ? _GEN_48 : _GEN_34; // @[elements.scala 123:26]
  wire  _GEN_53 = io_port_2_write_valid ? _GEN_49 : _GEN_35; // @[elements.scala 123:26]
  wire [64:0] _T_52 = {{1'd0}, io_port_3_read_in_bits_addr}; // @[elements.scala 118:104]
  wire [63:0] _T_56 = io_port_3_read_in_bits_addr + 64'h1; // @[elements.scala 118:104]
  wire  _GEN_55 = 2'h1 == _T_56[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_56 = 2'h2 == _T_56[1:0] ? content_2 : _GEN_55; // @[Cat.scala 29:58]
  wire  _GEN_57 = 2'h3 == _T_56[1:0] ? content_3 : _GEN_56; // @[Cat.scala 29:58]
  wire  _GEN_59 = 2'h1 == _T_52[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_60 = 2'h2 == _T_52[1:0] ? content_2 : _GEN_59; // @[Cat.scala 29:58]
  wire  _GEN_61 = 2'h3 == _T_52[1:0] ? content_3 : _GEN_60; // @[Cat.scala 29:58]
  wire [1:0] _T_58 = {_GEN_57,_GEN_61}; // @[Cat.scala 29:58]
  wire  _GEN_64 = 2'h0 == io_port_3_write_bits_addr[1:0] ? io_port_3_write_bits_value : _GEN_50; // @[elements.scala 124:49]
  wire  _GEN_65 = 2'h1 == io_port_3_write_bits_addr[1:0] ? io_port_3_write_bits_value : _GEN_51; // @[elements.scala 124:49]
  wire  _GEN_66 = 2'h2 == io_port_3_write_bits_addr[1:0] ? io_port_3_write_bits_value : _GEN_52; // @[elements.scala 124:49]
  wire  _GEN_67 = 2'h3 == io_port_3_write_bits_addr[1:0] ? io_port_3_write_bits_value : _GEN_53; // @[elements.scala 124:49]
  wire  _GEN_68 = io_port_3_write_valid ? _GEN_64 : _GEN_50; // @[elements.scala 123:26]
  wire  _GEN_69 = io_port_3_write_valid ? _GEN_65 : _GEN_51; // @[elements.scala 123:26]
  wire  _GEN_70 = io_port_3_write_valid ? _GEN_66 : _GEN_52; // @[elements.scala 123:26]
  wire  _GEN_71 = io_port_3_write_valid ? _GEN_67 : _GEN_53; // @[elements.scala 123:26]
  wire [64:0] _T_69 = {{1'd0}, io_port_4_read_in_bits_addr}; // @[elements.scala 118:104]
  wire [63:0] _T_73 = io_port_4_read_in_bits_addr + 64'h1; // @[elements.scala 118:104]
  wire  _GEN_73 = 2'h1 == _T_73[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_74 = 2'h2 == _T_73[1:0] ? content_2 : _GEN_73; // @[Cat.scala 29:58]
  wire  _GEN_75 = 2'h3 == _T_73[1:0] ? content_3 : _GEN_74; // @[Cat.scala 29:58]
  wire  _GEN_77 = 2'h1 == _T_69[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_78 = 2'h2 == _T_69[1:0] ? content_2 : _GEN_77; // @[Cat.scala 29:58]
  wire  _GEN_79 = 2'h3 == _T_69[1:0] ? content_3 : _GEN_78; // @[Cat.scala 29:58]
  wire [1:0] _T_75 = {_GEN_75,_GEN_79}; // @[Cat.scala 29:58]
  wire  _GEN_82 = 2'h0 == io_port_4_write_bits_addr[1:0] ? io_port_4_write_bits_value : _GEN_68; // @[elements.scala 124:49]
  wire  _GEN_83 = 2'h1 == io_port_4_write_bits_addr[1:0] ? io_port_4_write_bits_value : _GEN_69; // @[elements.scala 124:49]
  wire  _GEN_84 = 2'h2 == io_port_4_write_bits_addr[1:0] ? io_port_4_write_bits_value : _GEN_70; // @[elements.scala 124:49]
  wire  _GEN_85 = 2'h3 == io_port_4_write_bits_addr[1:0] ? io_port_4_write_bits_value : _GEN_71; // @[elements.scala 124:49]
  wire  _GEN_86 = io_port_4_write_valid ? _GEN_82 : _GEN_68; // @[elements.scala 123:26]
  wire  _GEN_87 = io_port_4_write_valid ? _GEN_83 : _GEN_69; // @[elements.scala 123:26]
  wire  _GEN_88 = io_port_4_write_valid ? _GEN_84 : _GEN_70; // @[elements.scala 123:26]
  wire  _GEN_89 = io_port_4_write_valid ? _GEN_85 : _GEN_71; // @[elements.scala 123:26]
  wire [64:0] _T_86 = {{1'd0}, io_port_5_read_in_bits_addr}; // @[elements.scala 118:104]
  wire [63:0] _T_90 = io_port_5_read_in_bits_addr + 64'h1; // @[elements.scala 118:104]
  wire  _GEN_91 = 2'h1 == _T_90[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_92 = 2'h2 == _T_90[1:0] ? content_2 : _GEN_91; // @[Cat.scala 29:58]
  wire  _GEN_93 = 2'h3 == _T_90[1:0] ? content_3 : _GEN_92; // @[Cat.scala 29:58]
  wire  _GEN_95 = 2'h1 == _T_86[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_96 = 2'h2 == _T_86[1:0] ? content_2 : _GEN_95; // @[Cat.scala 29:58]
  wire  _GEN_97 = 2'h3 == _T_86[1:0] ? content_3 : _GEN_96; // @[Cat.scala 29:58]
  wire [1:0] _T_92 = {_GEN_93,_GEN_97}; // @[Cat.scala 29:58]
  wire  _GEN_100 = 2'h0 == io_port_5_write_bits_addr[1:0] ? io_port_5_write_bits_value : _GEN_86; // @[elements.scala 124:49]
  wire  _GEN_101 = 2'h1 == io_port_5_write_bits_addr[1:0] ? io_port_5_write_bits_value : _GEN_87; // @[elements.scala 124:49]
  wire  _GEN_102 = 2'h2 == io_port_5_write_bits_addr[1:0] ? io_port_5_write_bits_value : _GEN_88; // @[elements.scala 124:49]
  wire  _GEN_103 = 2'h3 == io_port_5_write_bits_addr[1:0] ? io_port_5_write_bits_value : _GEN_89; // @[elements.scala 124:49]
  wire  _GEN_104 = io_port_5_write_valid ? _GEN_100 : _GEN_86; // @[elements.scala 123:26]
  wire  _GEN_105 = io_port_5_write_valid ? _GEN_101 : _GEN_87; // @[elements.scala 123:26]
  wire  _GEN_106 = io_port_5_write_valid ? _GEN_102 : _GEN_88; // @[elements.scala 123:26]
  wire  _GEN_107 = io_port_5_write_valid ? _GEN_103 : _GEN_89; // @[elements.scala 123:26]
  wire [64:0] _T_103 = {{1'd0}, io_port_6_read_in_bits_addr}; // @[elements.scala 118:104]
  wire [63:0] _T_107 = io_port_6_read_in_bits_addr + 64'h1; // @[elements.scala 118:104]
  wire  _GEN_109 = 2'h1 == _T_107[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_110 = 2'h2 == _T_107[1:0] ? content_2 : _GEN_109; // @[Cat.scala 29:58]
  wire  _GEN_111 = 2'h3 == _T_107[1:0] ? content_3 : _GEN_110; // @[Cat.scala 29:58]
  wire  _GEN_113 = 2'h1 == _T_103[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_114 = 2'h2 == _T_103[1:0] ? content_2 : _GEN_113; // @[Cat.scala 29:58]
  wire  _GEN_115 = 2'h3 == _T_103[1:0] ? content_3 : _GEN_114; // @[Cat.scala 29:58]
  wire [1:0] _T_109 = {_GEN_111,_GEN_115}; // @[Cat.scala 29:58]
  wire [64:0] _T_120 = {{1'd0}, io_port_7_read_in_bits_addr}; // @[elements.scala 118:104]
  wire [63:0] _T_124 = io_port_7_read_in_bits_addr + 64'h1; // @[elements.scala 118:104]
  wire  _GEN_127 = 2'h1 == _T_124[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_128 = 2'h2 == _T_124[1:0] ? content_2 : _GEN_127; // @[Cat.scala 29:58]
  wire  _GEN_129 = 2'h3 == _T_124[1:0] ? content_3 : _GEN_128; // @[Cat.scala 29:58]
  wire  _GEN_131 = 2'h1 == _T_120[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_132 = 2'h2 == _T_120[1:0] ? content_2 : _GEN_131; // @[Cat.scala 29:58]
  wire  _GEN_133 = 2'h3 == _T_120[1:0] ? content_3 : _GEN_132; // @[Cat.scala 29:58]
  wire [1:0] _T_126 = {_GEN_129,_GEN_133}; // @[Cat.scala 29:58]
  wire [64:0] _T_137 = {{1'd0}, io_port_8_read_in_bits_addr}; // @[elements.scala 118:104]
  wire [63:0] _T_141 = io_port_8_read_in_bits_addr + 64'h1; // @[elements.scala 118:104]
  wire  _GEN_145 = 2'h1 == _T_141[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_146 = 2'h2 == _T_141[1:0] ? content_2 : _GEN_145; // @[Cat.scala 29:58]
  wire  _GEN_147 = 2'h3 == _T_141[1:0] ? content_3 : _GEN_146; // @[Cat.scala 29:58]
  wire  _GEN_149 = 2'h1 == _T_137[1:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_150 = 2'h2 == _T_137[1:0] ? content_2 : _GEN_149; // @[Cat.scala 29:58]
  wire  _GEN_151 = 2'h3 == _T_137[1:0] ? content_3 : _GEN_150; // @[Cat.scala 29:58]
  wire [1:0] _T_143 = {_GEN_147,_GEN_151}; // @[Cat.scala 29:58]
  assign io_port_0_read_out_0 = io_port_0_read_in_valid & _T_7[0]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_0_read_out_1 = io_port_0_read_in_valid & _T_7[1]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_1_read_out_0 = io_port_1_read_in_valid & _T_24[0]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_1_read_out_1 = io_port_1_read_in_valid & _T_24[1]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_2_read_out_0 = io_port_2_read_in_valid & _T_41[0]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_2_read_out_1 = io_port_2_read_in_valid & _T_41[1]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_3_read_out_0 = io_port_3_read_in_valid & _T_58[0]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_3_read_out_1 = io_port_3_read_in_valid & _T_58[1]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_4_read_out_0 = io_port_4_read_in_valid & _T_75[0]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_4_read_out_1 = io_port_4_read_in_valid & _T_75[1]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_5_read_out_0 = io_port_5_read_in_valid & _T_92[0]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_5_read_out_1 = io_port_5_read_in_valid & _T_92[1]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_6_read_out_0 = io_port_6_read_in_valid & _T_109[0]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_6_read_out_1 = io_port_6_read_in_valid & _T_109[1]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_7_read_out_0 = io_port_7_read_in_valid & _T_126[0]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_7_read_out_1 = io_port_7_read_in_valid & _T_126[1]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_8_read_out_0 = io_port_8_read_in_valid & _T_143[0]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_8_read_out_1 = io_port_8_read_in_valid & _T_143[1]; // @[elements.scala 118:33 elements.scala 120:33]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  content_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  content_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  content_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  content_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      content_0 <= 1'h0;
    end else if (io_port_8_write_valid) begin
      if (2'h0 == io_port_8_write_bits_addr[1:0]) begin
        content_0 <= io_port_8_write_bits_value;
      end else if (io_port_7_write_valid) begin
        if (2'h0 == io_port_7_write_bits_addr[1:0]) begin
          content_0 <= io_port_7_write_bits_value;
        end else if (io_port_6_write_valid) begin
          if (2'h0 == io_port_6_write_bits_addr[1:0]) begin
            content_0 <= io_port_6_write_bits_value;
          end else if (io_port_5_write_valid) begin
            if (2'h0 == io_port_5_write_bits_addr[1:0]) begin
              content_0 <= io_port_5_write_bits_value;
            end else if (io_port_4_write_valid) begin
              if (2'h0 == io_port_4_write_bits_addr[1:0]) begin
                content_0 <= io_port_4_write_bits_value;
              end else if (io_port_3_write_valid) begin
                if (2'h0 == io_port_3_write_bits_addr[1:0]) begin
                  content_0 <= io_port_3_write_bits_value;
                end else if (io_port_2_write_valid) begin
                  if (2'h0 == io_port_2_write_bits_addr[1:0]) begin
                    content_0 <= io_port_2_write_bits_value;
                  end else if (io_port_1_write_valid) begin
                    if (2'h0 == io_port_1_write_bits_addr[1:0]) begin
                      content_0 <= io_port_1_write_bits_value;
                    end else if (io_port_0_write_valid) begin
                      if (2'h0 == io_port_0_write_bits_addr[1:0]) begin
                        content_0 <= io_port_0_write_bits_value;
                      end
                    end
                  end else if (io_port_0_write_valid) begin
                    if (2'h0 == io_port_0_write_bits_addr[1:0]) begin
                      content_0 <= io_port_0_write_bits_value;
                    end
                  end
                end else if (io_port_1_write_valid) begin
                  if (2'h0 == io_port_1_write_bits_addr[1:0]) begin
                    content_0 <= io_port_1_write_bits_value;
                  end else if (io_port_0_write_valid) begin
                    if (2'h0 == io_port_0_write_bits_addr[1:0]) begin
                      content_0 <= io_port_0_write_bits_value;
                    end
                  end
                end else if (io_port_0_write_valid) begin
                  if (2'h0 == io_port_0_write_bits_addr[1:0]) begin
                    content_0 <= io_port_0_write_bits_value;
                  end
                end
              end else if (io_port_2_write_valid) begin
                if (2'h0 == io_port_2_write_bits_addr[1:0]) begin
                  content_0 <= io_port_2_write_bits_value;
                end else if (io_port_1_write_valid) begin
                  if (2'h0 == io_port_1_write_bits_addr[1:0]) begin
                    content_0 <= io_port_1_write_bits_value;
                  end else begin
                    content_0 <= _GEN_14;
                  end
                end else begin
                  content_0 <= _GEN_14;
                end
              end else if (io_port_1_write_valid) begin
                if (2'h0 == io_port_1_write_bits_addr[1:0]) begin
                  content_0 <= io_port_1_write_bits_value;
                end else begin
                  content_0 <= _GEN_14;
                end
              end else begin
                content_0 <= _GEN_14;
              end
            end else if (io_port_3_write_valid) begin
              if (2'h0 == io_port_3_write_bits_addr[1:0]) begin
                content_0 <= io_port_3_write_bits_value;
              end else if (io_port_2_write_valid) begin
                if (2'h0 == io_port_2_write_bits_addr[1:0]) begin
                  content_0 <= io_port_2_write_bits_value;
                end else begin
                  content_0 <= _GEN_32;
                end
              end else begin
                content_0 <= _GEN_32;
              end
            end else if (io_port_2_write_valid) begin
              if (2'h0 == io_port_2_write_bits_addr[1:0]) begin
                content_0 <= io_port_2_write_bits_value;
              end else begin
                content_0 <= _GEN_32;
              end
            end else begin
              content_0 <= _GEN_32;
            end
          end else if (io_port_4_write_valid) begin
            if (2'h0 == io_port_4_write_bits_addr[1:0]) begin
              content_0 <= io_port_4_write_bits_value;
            end else if (io_port_3_write_valid) begin
              if (2'h0 == io_port_3_write_bits_addr[1:0]) begin
                content_0 <= io_port_3_write_bits_value;
              end else begin
                content_0 <= _GEN_50;
              end
            end else begin
              content_0 <= _GEN_50;
            end
          end else if (io_port_3_write_valid) begin
            if (2'h0 == io_port_3_write_bits_addr[1:0]) begin
              content_0 <= io_port_3_write_bits_value;
            end else begin
              content_0 <= _GEN_50;
            end
          end else begin
            content_0 <= _GEN_50;
          end
        end else if (io_port_5_write_valid) begin
          if (2'h0 == io_port_5_write_bits_addr[1:0]) begin
            content_0 <= io_port_5_write_bits_value;
          end else if (io_port_4_write_valid) begin
            if (2'h0 == io_port_4_write_bits_addr[1:0]) begin
              content_0 <= io_port_4_write_bits_value;
            end else begin
              content_0 <= _GEN_68;
            end
          end else begin
            content_0 <= _GEN_68;
          end
        end else if (io_port_4_write_valid) begin
          if (2'h0 == io_port_4_write_bits_addr[1:0]) begin
            content_0 <= io_port_4_write_bits_value;
          end else begin
            content_0 <= _GEN_68;
          end
        end else begin
          content_0 <= _GEN_68;
        end
      end else if (io_port_6_write_valid) begin
        if (2'h0 == io_port_6_write_bits_addr[1:0]) begin
          content_0 <= io_port_6_write_bits_value;
        end else if (io_port_5_write_valid) begin
          if (2'h0 == io_port_5_write_bits_addr[1:0]) begin
            content_0 <= io_port_5_write_bits_value;
          end else begin
            content_0 <= _GEN_86;
          end
        end else begin
          content_0 <= _GEN_86;
        end
      end else if (io_port_5_write_valid) begin
        if (2'h0 == io_port_5_write_bits_addr[1:0]) begin
          content_0 <= io_port_5_write_bits_value;
        end else begin
          content_0 <= _GEN_86;
        end
      end else begin
        content_0 <= _GEN_86;
      end
    end else if (io_port_7_write_valid) begin
      if (2'h0 == io_port_7_write_bits_addr[1:0]) begin
        content_0 <= io_port_7_write_bits_value;
      end else if (io_port_6_write_valid) begin
        if (2'h0 == io_port_6_write_bits_addr[1:0]) begin
          content_0 <= io_port_6_write_bits_value;
        end else begin
          content_0 <= _GEN_104;
        end
      end else begin
        content_0 <= _GEN_104;
      end
    end else if (io_port_6_write_valid) begin
      if (2'h0 == io_port_6_write_bits_addr[1:0]) begin
        content_0 <= io_port_6_write_bits_value;
      end else begin
        content_0 <= _GEN_104;
      end
    end else begin
      content_0 <= _GEN_104;
    end
    if (reset) begin
      content_1 <= 1'h0;
    end else if (io_port_8_write_valid) begin
      if (2'h1 == io_port_8_write_bits_addr[1:0]) begin
        content_1 <= io_port_8_write_bits_value;
      end else if (io_port_7_write_valid) begin
        if (2'h1 == io_port_7_write_bits_addr[1:0]) begin
          content_1 <= io_port_7_write_bits_value;
        end else if (io_port_6_write_valid) begin
          if (2'h1 == io_port_6_write_bits_addr[1:0]) begin
            content_1 <= io_port_6_write_bits_value;
          end else if (io_port_5_write_valid) begin
            if (2'h1 == io_port_5_write_bits_addr[1:0]) begin
              content_1 <= io_port_5_write_bits_value;
            end else if (io_port_4_write_valid) begin
              if (2'h1 == io_port_4_write_bits_addr[1:0]) begin
                content_1 <= io_port_4_write_bits_value;
              end else if (io_port_3_write_valid) begin
                if (2'h1 == io_port_3_write_bits_addr[1:0]) begin
                  content_1 <= io_port_3_write_bits_value;
                end else if (io_port_2_write_valid) begin
                  if (2'h1 == io_port_2_write_bits_addr[1:0]) begin
                    content_1 <= io_port_2_write_bits_value;
                  end else if (io_port_1_write_valid) begin
                    if (2'h1 == io_port_1_write_bits_addr[1:0]) begin
                      content_1 <= io_port_1_write_bits_value;
                    end else if (io_port_0_write_valid) begin
                      if (2'h1 == io_port_0_write_bits_addr[1:0]) begin
                        content_1 <= io_port_0_write_bits_value;
                      end
                    end
                  end else if (io_port_0_write_valid) begin
                    if (2'h1 == io_port_0_write_bits_addr[1:0]) begin
                      content_1 <= io_port_0_write_bits_value;
                    end
                  end
                end else if (io_port_1_write_valid) begin
                  if (2'h1 == io_port_1_write_bits_addr[1:0]) begin
                    content_1 <= io_port_1_write_bits_value;
                  end else if (io_port_0_write_valid) begin
                    if (2'h1 == io_port_0_write_bits_addr[1:0]) begin
                      content_1 <= io_port_0_write_bits_value;
                    end
                  end
                end else if (io_port_0_write_valid) begin
                  if (2'h1 == io_port_0_write_bits_addr[1:0]) begin
                    content_1 <= io_port_0_write_bits_value;
                  end
                end
              end else if (io_port_2_write_valid) begin
                if (2'h1 == io_port_2_write_bits_addr[1:0]) begin
                  content_1 <= io_port_2_write_bits_value;
                end else if (io_port_1_write_valid) begin
                  if (2'h1 == io_port_1_write_bits_addr[1:0]) begin
                    content_1 <= io_port_1_write_bits_value;
                  end else begin
                    content_1 <= _GEN_15;
                  end
                end else begin
                  content_1 <= _GEN_15;
                end
              end else if (io_port_1_write_valid) begin
                if (2'h1 == io_port_1_write_bits_addr[1:0]) begin
                  content_1 <= io_port_1_write_bits_value;
                end else begin
                  content_1 <= _GEN_15;
                end
              end else begin
                content_1 <= _GEN_15;
              end
            end else if (io_port_3_write_valid) begin
              if (2'h1 == io_port_3_write_bits_addr[1:0]) begin
                content_1 <= io_port_3_write_bits_value;
              end else if (io_port_2_write_valid) begin
                if (2'h1 == io_port_2_write_bits_addr[1:0]) begin
                  content_1 <= io_port_2_write_bits_value;
                end else begin
                  content_1 <= _GEN_33;
                end
              end else begin
                content_1 <= _GEN_33;
              end
            end else if (io_port_2_write_valid) begin
              if (2'h1 == io_port_2_write_bits_addr[1:0]) begin
                content_1 <= io_port_2_write_bits_value;
              end else begin
                content_1 <= _GEN_33;
              end
            end else begin
              content_1 <= _GEN_33;
            end
          end else if (io_port_4_write_valid) begin
            if (2'h1 == io_port_4_write_bits_addr[1:0]) begin
              content_1 <= io_port_4_write_bits_value;
            end else if (io_port_3_write_valid) begin
              if (2'h1 == io_port_3_write_bits_addr[1:0]) begin
                content_1 <= io_port_3_write_bits_value;
              end else begin
                content_1 <= _GEN_51;
              end
            end else begin
              content_1 <= _GEN_51;
            end
          end else if (io_port_3_write_valid) begin
            if (2'h1 == io_port_3_write_bits_addr[1:0]) begin
              content_1 <= io_port_3_write_bits_value;
            end else begin
              content_1 <= _GEN_51;
            end
          end else begin
            content_1 <= _GEN_51;
          end
        end else if (io_port_5_write_valid) begin
          if (2'h1 == io_port_5_write_bits_addr[1:0]) begin
            content_1 <= io_port_5_write_bits_value;
          end else if (io_port_4_write_valid) begin
            if (2'h1 == io_port_4_write_bits_addr[1:0]) begin
              content_1 <= io_port_4_write_bits_value;
            end else begin
              content_1 <= _GEN_69;
            end
          end else begin
            content_1 <= _GEN_69;
          end
        end else if (io_port_4_write_valid) begin
          if (2'h1 == io_port_4_write_bits_addr[1:0]) begin
            content_1 <= io_port_4_write_bits_value;
          end else begin
            content_1 <= _GEN_69;
          end
        end else begin
          content_1 <= _GEN_69;
        end
      end else if (io_port_6_write_valid) begin
        if (2'h1 == io_port_6_write_bits_addr[1:0]) begin
          content_1 <= io_port_6_write_bits_value;
        end else if (io_port_5_write_valid) begin
          if (2'h1 == io_port_5_write_bits_addr[1:0]) begin
            content_1 <= io_port_5_write_bits_value;
          end else begin
            content_1 <= _GEN_87;
          end
        end else begin
          content_1 <= _GEN_87;
        end
      end else if (io_port_5_write_valid) begin
        if (2'h1 == io_port_5_write_bits_addr[1:0]) begin
          content_1 <= io_port_5_write_bits_value;
        end else begin
          content_1 <= _GEN_87;
        end
      end else begin
        content_1 <= _GEN_87;
      end
    end else if (io_port_7_write_valid) begin
      if (2'h1 == io_port_7_write_bits_addr[1:0]) begin
        content_1 <= io_port_7_write_bits_value;
      end else if (io_port_6_write_valid) begin
        if (2'h1 == io_port_6_write_bits_addr[1:0]) begin
          content_1 <= io_port_6_write_bits_value;
        end else begin
          content_1 <= _GEN_105;
        end
      end else begin
        content_1 <= _GEN_105;
      end
    end else if (io_port_6_write_valid) begin
      if (2'h1 == io_port_6_write_bits_addr[1:0]) begin
        content_1 <= io_port_6_write_bits_value;
      end else begin
        content_1 <= _GEN_105;
      end
    end else begin
      content_1 <= _GEN_105;
    end
    if (reset) begin
      content_2 <= 1'h0;
    end else if (io_port_8_write_valid) begin
      if (2'h2 == io_port_8_write_bits_addr[1:0]) begin
        content_2 <= io_port_8_write_bits_value;
      end else if (io_port_7_write_valid) begin
        if (2'h2 == io_port_7_write_bits_addr[1:0]) begin
          content_2 <= io_port_7_write_bits_value;
        end else if (io_port_6_write_valid) begin
          if (2'h2 == io_port_6_write_bits_addr[1:0]) begin
            content_2 <= io_port_6_write_bits_value;
          end else if (io_port_5_write_valid) begin
            if (2'h2 == io_port_5_write_bits_addr[1:0]) begin
              content_2 <= io_port_5_write_bits_value;
            end else if (io_port_4_write_valid) begin
              if (2'h2 == io_port_4_write_bits_addr[1:0]) begin
                content_2 <= io_port_4_write_bits_value;
              end else if (io_port_3_write_valid) begin
                if (2'h2 == io_port_3_write_bits_addr[1:0]) begin
                  content_2 <= io_port_3_write_bits_value;
                end else if (io_port_2_write_valid) begin
                  if (2'h2 == io_port_2_write_bits_addr[1:0]) begin
                    content_2 <= io_port_2_write_bits_value;
                  end else if (io_port_1_write_valid) begin
                    if (2'h2 == io_port_1_write_bits_addr[1:0]) begin
                      content_2 <= io_port_1_write_bits_value;
                    end else if (io_port_0_write_valid) begin
                      if (2'h2 == io_port_0_write_bits_addr[1:0]) begin
                        content_2 <= io_port_0_write_bits_value;
                      end
                    end
                  end else if (io_port_0_write_valid) begin
                    if (2'h2 == io_port_0_write_bits_addr[1:0]) begin
                      content_2 <= io_port_0_write_bits_value;
                    end
                  end
                end else if (io_port_1_write_valid) begin
                  if (2'h2 == io_port_1_write_bits_addr[1:0]) begin
                    content_2 <= io_port_1_write_bits_value;
                  end else if (io_port_0_write_valid) begin
                    if (2'h2 == io_port_0_write_bits_addr[1:0]) begin
                      content_2 <= io_port_0_write_bits_value;
                    end
                  end
                end else if (io_port_0_write_valid) begin
                  if (2'h2 == io_port_0_write_bits_addr[1:0]) begin
                    content_2 <= io_port_0_write_bits_value;
                  end
                end
              end else if (io_port_2_write_valid) begin
                if (2'h2 == io_port_2_write_bits_addr[1:0]) begin
                  content_2 <= io_port_2_write_bits_value;
                end else if (io_port_1_write_valid) begin
                  if (2'h2 == io_port_1_write_bits_addr[1:0]) begin
                    content_2 <= io_port_1_write_bits_value;
                  end else begin
                    content_2 <= _GEN_16;
                  end
                end else begin
                  content_2 <= _GEN_16;
                end
              end else if (io_port_1_write_valid) begin
                if (2'h2 == io_port_1_write_bits_addr[1:0]) begin
                  content_2 <= io_port_1_write_bits_value;
                end else begin
                  content_2 <= _GEN_16;
                end
              end else begin
                content_2 <= _GEN_16;
              end
            end else if (io_port_3_write_valid) begin
              if (2'h2 == io_port_3_write_bits_addr[1:0]) begin
                content_2 <= io_port_3_write_bits_value;
              end else if (io_port_2_write_valid) begin
                if (2'h2 == io_port_2_write_bits_addr[1:0]) begin
                  content_2 <= io_port_2_write_bits_value;
                end else begin
                  content_2 <= _GEN_34;
                end
              end else begin
                content_2 <= _GEN_34;
              end
            end else if (io_port_2_write_valid) begin
              if (2'h2 == io_port_2_write_bits_addr[1:0]) begin
                content_2 <= io_port_2_write_bits_value;
              end else begin
                content_2 <= _GEN_34;
              end
            end else begin
              content_2 <= _GEN_34;
            end
          end else if (io_port_4_write_valid) begin
            if (2'h2 == io_port_4_write_bits_addr[1:0]) begin
              content_2 <= io_port_4_write_bits_value;
            end else if (io_port_3_write_valid) begin
              if (2'h2 == io_port_3_write_bits_addr[1:0]) begin
                content_2 <= io_port_3_write_bits_value;
              end else begin
                content_2 <= _GEN_52;
              end
            end else begin
              content_2 <= _GEN_52;
            end
          end else if (io_port_3_write_valid) begin
            if (2'h2 == io_port_3_write_bits_addr[1:0]) begin
              content_2 <= io_port_3_write_bits_value;
            end else begin
              content_2 <= _GEN_52;
            end
          end else begin
            content_2 <= _GEN_52;
          end
        end else if (io_port_5_write_valid) begin
          if (2'h2 == io_port_5_write_bits_addr[1:0]) begin
            content_2 <= io_port_5_write_bits_value;
          end else if (io_port_4_write_valid) begin
            if (2'h2 == io_port_4_write_bits_addr[1:0]) begin
              content_2 <= io_port_4_write_bits_value;
            end else begin
              content_2 <= _GEN_70;
            end
          end else begin
            content_2 <= _GEN_70;
          end
        end else if (io_port_4_write_valid) begin
          if (2'h2 == io_port_4_write_bits_addr[1:0]) begin
            content_2 <= io_port_4_write_bits_value;
          end else begin
            content_2 <= _GEN_70;
          end
        end else begin
          content_2 <= _GEN_70;
        end
      end else if (io_port_6_write_valid) begin
        if (2'h2 == io_port_6_write_bits_addr[1:0]) begin
          content_2 <= io_port_6_write_bits_value;
        end else if (io_port_5_write_valid) begin
          if (2'h2 == io_port_5_write_bits_addr[1:0]) begin
            content_2 <= io_port_5_write_bits_value;
          end else begin
            content_2 <= _GEN_88;
          end
        end else begin
          content_2 <= _GEN_88;
        end
      end else if (io_port_5_write_valid) begin
        if (2'h2 == io_port_5_write_bits_addr[1:0]) begin
          content_2 <= io_port_5_write_bits_value;
        end else begin
          content_2 <= _GEN_88;
        end
      end else begin
        content_2 <= _GEN_88;
      end
    end else if (io_port_7_write_valid) begin
      if (2'h2 == io_port_7_write_bits_addr[1:0]) begin
        content_2 <= io_port_7_write_bits_value;
      end else if (io_port_6_write_valid) begin
        if (2'h2 == io_port_6_write_bits_addr[1:0]) begin
          content_2 <= io_port_6_write_bits_value;
        end else begin
          content_2 <= _GEN_106;
        end
      end else begin
        content_2 <= _GEN_106;
      end
    end else if (io_port_6_write_valid) begin
      if (2'h2 == io_port_6_write_bits_addr[1:0]) begin
        content_2 <= io_port_6_write_bits_value;
      end else begin
        content_2 <= _GEN_106;
      end
    end else begin
      content_2 <= _GEN_106;
    end
    if (reset) begin
      content_3 <= 1'h0;
    end else if (io_port_8_write_valid) begin
      if (2'h3 == io_port_8_write_bits_addr[1:0]) begin
        content_3 <= io_port_8_write_bits_value;
      end else if (io_port_7_write_valid) begin
        if (2'h3 == io_port_7_write_bits_addr[1:0]) begin
          content_3 <= io_port_7_write_bits_value;
        end else if (io_port_6_write_valid) begin
          if (2'h3 == io_port_6_write_bits_addr[1:0]) begin
            content_3 <= io_port_6_write_bits_value;
          end else if (io_port_5_write_valid) begin
            if (2'h3 == io_port_5_write_bits_addr[1:0]) begin
              content_3 <= io_port_5_write_bits_value;
            end else if (io_port_4_write_valid) begin
              if (2'h3 == io_port_4_write_bits_addr[1:0]) begin
                content_3 <= io_port_4_write_bits_value;
              end else if (io_port_3_write_valid) begin
                if (2'h3 == io_port_3_write_bits_addr[1:0]) begin
                  content_3 <= io_port_3_write_bits_value;
                end else if (io_port_2_write_valid) begin
                  if (2'h3 == io_port_2_write_bits_addr[1:0]) begin
                    content_3 <= io_port_2_write_bits_value;
                  end else if (io_port_1_write_valid) begin
                    if (2'h3 == io_port_1_write_bits_addr[1:0]) begin
                      content_3 <= io_port_1_write_bits_value;
                    end else if (io_port_0_write_valid) begin
                      if (2'h3 == io_port_0_write_bits_addr[1:0]) begin
                        content_3 <= io_port_0_write_bits_value;
                      end
                    end
                  end else if (io_port_0_write_valid) begin
                    if (2'h3 == io_port_0_write_bits_addr[1:0]) begin
                      content_3 <= io_port_0_write_bits_value;
                    end
                  end
                end else if (io_port_1_write_valid) begin
                  if (2'h3 == io_port_1_write_bits_addr[1:0]) begin
                    content_3 <= io_port_1_write_bits_value;
                  end else if (io_port_0_write_valid) begin
                    if (2'h3 == io_port_0_write_bits_addr[1:0]) begin
                      content_3 <= io_port_0_write_bits_value;
                    end
                  end
                end else if (io_port_0_write_valid) begin
                  if (2'h3 == io_port_0_write_bits_addr[1:0]) begin
                    content_3 <= io_port_0_write_bits_value;
                  end
                end
              end else if (io_port_2_write_valid) begin
                if (2'h3 == io_port_2_write_bits_addr[1:0]) begin
                  content_3 <= io_port_2_write_bits_value;
                end else if (io_port_1_write_valid) begin
                  if (2'h3 == io_port_1_write_bits_addr[1:0]) begin
                    content_3 <= io_port_1_write_bits_value;
                  end else begin
                    content_3 <= _GEN_17;
                  end
                end else begin
                  content_3 <= _GEN_17;
                end
              end else if (io_port_1_write_valid) begin
                if (2'h3 == io_port_1_write_bits_addr[1:0]) begin
                  content_3 <= io_port_1_write_bits_value;
                end else begin
                  content_3 <= _GEN_17;
                end
              end else begin
                content_3 <= _GEN_17;
              end
            end else if (io_port_3_write_valid) begin
              if (2'h3 == io_port_3_write_bits_addr[1:0]) begin
                content_3 <= io_port_3_write_bits_value;
              end else if (io_port_2_write_valid) begin
                if (2'h3 == io_port_2_write_bits_addr[1:0]) begin
                  content_3 <= io_port_2_write_bits_value;
                end else begin
                  content_3 <= _GEN_35;
                end
              end else begin
                content_3 <= _GEN_35;
              end
            end else if (io_port_2_write_valid) begin
              if (2'h3 == io_port_2_write_bits_addr[1:0]) begin
                content_3 <= io_port_2_write_bits_value;
              end else begin
                content_3 <= _GEN_35;
              end
            end else begin
              content_3 <= _GEN_35;
            end
          end else if (io_port_4_write_valid) begin
            if (2'h3 == io_port_4_write_bits_addr[1:0]) begin
              content_3 <= io_port_4_write_bits_value;
            end else if (io_port_3_write_valid) begin
              if (2'h3 == io_port_3_write_bits_addr[1:0]) begin
                content_3 <= io_port_3_write_bits_value;
              end else begin
                content_3 <= _GEN_53;
              end
            end else begin
              content_3 <= _GEN_53;
            end
          end else if (io_port_3_write_valid) begin
            if (2'h3 == io_port_3_write_bits_addr[1:0]) begin
              content_3 <= io_port_3_write_bits_value;
            end else begin
              content_3 <= _GEN_53;
            end
          end else begin
            content_3 <= _GEN_53;
          end
        end else if (io_port_5_write_valid) begin
          if (2'h3 == io_port_5_write_bits_addr[1:0]) begin
            content_3 <= io_port_5_write_bits_value;
          end else if (io_port_4_write_valid) begin
            if (2'h3 == io_port_4_write_bits_addr[1:0]) begin
              content_3 <= io_port_4_write_bits_value;
            end else begin
              content_3 <= _GEN_71;
            end
          end else begin
            content_3 <= _GEN_71;
          end
        end else if (io_port_4_write_valid) begin
          if (2'h3 == io_port_4_write_bits_addr[1:0]) begin
            content_3 <= io_port_4_write_bits_value;
          end else begin
            content_3 <= _GEN_71;
          end
        end else begin
          content_3 <= _GEN_71;
        end
      end else if (io_port_6_write_valid) begin
        if (2'h3 == io_port_6_write_bits_addr[1:0]) begin
          content_3 <= io_port_6_write_bits_value;
        end else if (io_port_5_write_valid) begin
          if (2'h3 == io_port_5_write_bits_addr[1:0]) begin
            content_3 <= io_port_5_write_bits_value;
          end else begin
            content_3 <= _GEN_89;
          end
        end else begin
          content_3 <= _GEN_89;
        end
      end else if (io_port_5_write_valid) begin
        if (2'h3 == io_port_5_write_bits_addr[1:0]) begin
          content_3 <= io_port_5_write_bits_value;
        end else begin
          content_3 <= _GEN_89;
        end
      end else begin
        content_3 <= _GEN_89;
      end
    end else if (io_port_7_write_valid) begin
      if (2'h3 == io_port_7_write_bits_addr[1:0]) begin
        content_3 <= io_port_7_write_bits_value;
      end else if (io_port_6_write_valid) begin
        if (2'h3 == io_port_6_write_bits_addr[1:0]) begin
          content_3 <= io_port_6_write_bits_value;
        end else begin
          content_3 <= _GEN_107;
        end
      end else begin
        content_3 <= _GEN_107;
      end
    end else if (io_port_6_write_valid) begin
      if (2'h3 == io_port_6_write_bits_addr[1:0]) begin
        content_3 <= io_port_6_write_bits_value;
      end else begin
        content_3 <= _GEN_107;
      end
    end else begin
      content_3 <= _GEN_107;
    end
  end
endmodule
module Arbiter_2(
  input         io_in_0_valid,
  input  [1:0]  io_in_0_bits_bank,
  input         io_in_0_bits_address,
  input  [30:0] io_in_0_bits_inputValue_0_tag,
  input  [30:0] io_in_0_bits_inputValue_1_tag,
  input         io_in_1_valid,
  input  [1:0]  io_in_1_bits_bank,
  input         io_in_1_bits_address,
  input  [30:0] io_in_1_bits_inputValue_0_tag,
  input  [30:0] io_in_1_bits_inputValue_1_tag,
  input         io_in_2_valid,
  input  [1:0]  io_in_2_bits_bank,
  input         io_in_2_bits_address,
  input  [30:0] io_in_2_bits_inputValue_0_tag,
  input  [30:0] io_in_2_bits_inputValue_1_tag,
  input         io_in_3_valid,
  input  [1:0]  io_in_3_bits_bank,
  input         io_in_3_bits_address,
  input  [30:0] io_in_3_bits_inputValue_0_tag,
  input  [30:0] io_in_3_bits_inputValue_1_tag,
  input         io_in_4_valid,
  input  [1:0]  io_in_4_bits_bank,
  input         io_in_4_bits_address,
  input  [30:0] io_in_4_bits_inputValue_0_tag,
  input  [30:0] io_in_4_bits_inputValue_1_tag,
  input         io_in_5_valid,
  input  [1:0]  io_in_5_bits_bank,
  input         io_in_5_bits_address,
  input  [30:0] io_in_5_bits_inputValue_0_tag,
  input  [30:0] io_in_5_bits_inputValue_1_tag,
  input         io_in_6_valid,
  input  [1:0]  io_in_6_bits_bank,
  input         io_in_6_bits_address,
  input  [30:0] io_in_6_bits_inputValue_0_tag,
  input  [30:0] io_in_6_bits_inputValue_1_tag,
  input         io_in_7_valid,
  input  [1:0]  io_in_7_bits_bank,
  input         io_in_7_bits_address,
  input  [30:0] io_in_7_bits_inputValue_0_tag,
  input  [30:0] io_in_7_bits_inputValue_1_tag,
  output        io_out_valid,
  output [1:0]  io_out_bits_bank,
  output        io_out_bits_address,
  output [30:0] io_out_bits_inputValue_0_tag,
  output [30:0] io_out_bits_inputValue_1_tag
);
  wire [30:0] _GEN_1 = io_in_6_valid ? io_in_6_bits_inputValue_0_tag : io_in_7_bits_inputValue_0_tag; // @[Arbiter.scala 126:27]
  wire [30:0] _GEN_2 = io_in_6_valid ? io_in_6_bits_inputValue_1_tag : io_in_7_bits_inputValue_1_tag; // @[Arbiter.scala 126:27]
  wire  _GEN_3 = io_in_6_valid ? io_in_6_bits_address : io_in_7_bits_address; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_4 = io_in_6_valid ? io_in_6_bits_bank : io_in_7_bits_bank; // @[Arbiter.scala 126:27]
  wire [30:0] _GEN_6 = io_in_5_valid ? io_in_5_bits_inputValue_0_tag : _GEN_1; // @[Arbiter.scala 126:27]
  wire [30:0] _GEN_7 = io_in_5_valid ? io_in_5_bits_inputValue_1_tag : _GEN_2; // @[Arbiter.scala 126:27]
  wire  _GEN_8 = io_in_5_valid ? io_in_5_bits_address : _GEN_3; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_9 = io_in_5_valid ? io_in_5_bits_bank : _GEN_4; // @[Arbiter.scala 126:27]
  wire [30:0] _GEN_11 = io_in_4_valid ? io_in_4_bits_inputValue_0_tag : _GEN_6; // @[Arbiter.scala 126:27]
  wire [30:0] _GEN_12 = io_in_4_valid ? io_in_4_bits_inputValue_1_tag : _GEN_7; // @[Arbiter.scala 126:27]
  wire  _GEN_13 = io_in_4_valid ? io_in_4_bits_address : _GEN_8; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_14 = io_in_4_valid ? io_in_4_bits_bank : _GEN_9; // @[Arbiter.scala 126:27]
  wire [30:0] _GEN_16 = io_in_3_valid ? io_in_3_bits_inputValue_0_tag : _GEN_11; // @[Arbiter.scala 126:27]
  wire [30:0] _GEN_17 = io_in_3_valid ? io_in_3_bits_inputValue_1_tag : _GEN_12; // @[Arbiter.scala 126:27]
  wire  _GEN_18 = io_in_3_valid ? io_in_3_bits_address : _GEN_13; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_19 = io_in_3_valid ? io_in_3_bits_bank : _GEN_14; // @[Arbiter.scala 126:27]
  wire [30:0] _GEN_21 = io_in_2_valid ? io_in_2_bits_inputValue_0_tag : _GEN_16; // @[Arbiter.scala 126:27]
  wire [30:0] _GEN_22 = io_in_2_valid ? io_in_2_bits_inputValue_1_tag : _GEN_17; // @[Arbiter.scala 126:27]
  wire  _GEN_23 = io_in_2_valid ? io_in_2_bits_address : _GEN_18; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_24 = io_in_2_valid ? io_in_2_bits_bank : _GEN_19; // @[Arbiter.scala 126:27]
  wire [30:0] _GEN_26 = io_in_1_valid ? io_in_1_bits_inputValue_0_tag : _GEN_21; // @[Arbiter.scala 126:27]
  wire [30:0] _GEN_27 = io_in_1_valid ? io_in_1_bits_inputValue_1_tag : _GEN_22; // @[Arbiter.scala 126:27]
  wire  _GEN_28 = io_in_1_valid ? io_in_1_bits_address : _GEN_23; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_29 = io_in_1_valid ? io_in_1_bits_bank : _GEN_24; // @[Arbiter.scala 126:27]
  wire  _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  _T_1 = _T | io_in_2_valid; // @[Arbiter.scala 31:68]
  wire  _T_2 = _T_1 | io_in_3_valid; // @[Arbiter.scala 31:68]
  wire  _T_3 = _T_2 | io_in_4_valid; // @[Arbiter.scala 31:68]
  wire  _T_4 = _T_3 | io_in_5_valid; // @[Arbiter.scala 31:68]
  wire  _T_5 = _T_4 | io_in_6_valid; // @[Arbiter.scala 31:68]
  wire  grant_7 = ~_T_5; // @[Arbiter.scala 31:78]
  wire  _T_14 = ~grant_7; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_14 | io_in_7_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_bank = io_in_0_valid ? io_in_0_bits_bank : _GEN_29; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_address = io_in_0_valid ? io_in_0_bits_address : _GEN_28; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_inputValue_0_tag = io_in_0_valid ? io_in_0_bits_inputValue_0_tag : _GEN_26; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_inputValue_1_tag = io_in_0_valid ? io_in_0_bits_inputValue_1_tag : _GEN_27; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
endmodule
module Gem5Cache(
  input         clock,
  input         reset,
  input         io_cpu_0_req_valid,
  input  [31:0] io_cpu_0_req_bits_addr,
  input  [27:0] io_cpu_0_req_bits_command,
  input  [1:0]  io_cpu_0_req_bits_way,
  input  [1:0]  io_cpu_0_req_bits_replaceWay,
  output        io_cpu_0_resp_valid,
  output        io_cpu_0_resp_bits_iswrite,
  output [1:0]  io_cpu_0_resp_bits_way,
  input         io_cpu_1_req_valid,
  input  [31:0] io_cpu_1_req_bits_addr,
  input  [27:0] io_cpu_1_req_bits_command,
  input  [1:0]  io_cpu_1_req_bits_way,
  input  [1:0]  io_cpu_1_req_bits_replaceWay,
  output        io_cpu_1_resp_valid,
  output        io_cpu_1_resp_bits_iswrite,
  output [1:0]  io_cpu_1_resp_bits_way,
  input         io_cpu_2_req_valid,
  input  [31:0] io_cpu_2_req_bits_addr,
  input  [27:0] io_cpu_2_req_bits_command,
  input  [1:0]  io_cpu_2_req_bits_way,
  input  [1:0]  io_cpu_2_req_bits_replaceWay,
  output        io_cpu_2_resp_valid,
  output        io_cpu_2_resp_bits_iswrite,
  output [1:0]  io_cpu_2_resp_bits_way,
  input         io_cpu_3_req_valid,
  input  [31:0] io_cpu_3_req_bits_addr,
  input  [27:0] io_cpu_3_req_bits_command,
  input  [1:0]  io_cpu_3_req_bits_way,
  input  [1:0]  io_cpu_3_req_bits_replaceWay,
  output        io_cpu_3_resp_valid,
  output        io_cpu_3_resp_bits_iswrite,
  output [1:0]  io_cpu_3_resp_bits_way,
  input         io_cpu_4_req_valid,
  input  [31:0] io_cpu_4_req_bits_addr,
  input  [27:0] io_cpu_4_req_bits_command,
  input  [1:0]  io_cpu_4_req_bits_way,
  input  [1:0]  io_cpu_4_req_bits_replaceWay,
  output        io_cpu_4_resp_valid,
  output        io_cpu_4_resp_bits_iswrite,
  output [1:0]  io_cpu_4_resp_bits_way,
  input         io_cpu_5_req_valid,
  input  [31:0] io_cpu_5_req_bits_addr,
  input  [27:0] io_cpu_5_req_bits_command,
  input  [1:0]  io_cpu_5_req_bits_way,
  input  [1:0]  io_cpu_5_req_bits_replaceWay,
  output        io_cpu_5_resp_valid,
  output        io_cpu_5_resp_bits_iswrite,
  output [1:0]  io_cpu_5_resp_bits_way,
  input         io_cpu_6_req_valid,
  input  [31:0] io_cpu_6_req_bits_addr,
  input  [27:0] io_cpu_6_req_bits_command,
  input  [1:0]  io_cpu_6_req_bits_way,
  input  [1:0]  io_cpu_6_req_bits_replaceWay,
  output        io_cpu_6_resp_valid,
  output        io_cpu_6_resp_bits_iswrite,
  output [1:0]  io_cpu_6_resp_bits_way,
  input         io_cpu_7_req_valid,
  input  [31:0] io_cpu_7_req_bits_addr,
  input  [63:0] io_cpu_7_req_bits_data,
  input  [27:0] io_cpu_7_req_bits_command,
  input  [1:0]  io_cpu_7_req_bits_way,
  input  [1:0]  io_cpu_7_req_bits_replaceWay,
  output        io_cpu_7_resp_valid,
  output        io_cpu_7_resp_bits_iswrite,
  output [1:0]  io_cpu_7_resp_bits_way,
  input         io_probe_req_valid,
  input  [31:0] io_probe_req_bits_addr,
  input  [27:0] io_probe_req_bits_command,
  output        io_probe_resp_valid,
  output [1:0]  io_probe_resp_bits_way,
  output        io_probe_multiWay_valid,
  output [1:0]  io_probe_multiWay_bits_way_0,
  output [1:0]  io_probe_multiWay_bits_way_1,
  output [31:0] io_probe_multiWay_bits_addr,
  input         io_bipassLD_in_valid,
  input  [31:0] io_bipassLD_in_bits_addr,
  input  [2:0]  io_bipassLD_in_bits_way,
  output        io_bipassLD_out_valid,
  output [63:0] io_bipassLD_out_bits_data
);
  wire  biPassModule_clock; // @[AXICache.scala 61:28]
  wire  biPassModule_reset; // @[AXICache.scala 61:28]
  wire  biPassModule_io_in_valid; // @[AXICache.scala 61:28]
  wire [31:0] biPassModule_io_in_bits_addr; // @[AXICache.scala 61:28]
  wire [2:0] biPassModule_io_in_bits_way; // @[AXICache.scala 61:28]
  wire  biPassModule_io_dataMem_in_valid; // @[AXICache.scala 61:28]
  wire [31:0] biPassModule_io_dataMem_in_bits_address; // @[AXICache.scala 61:28]
  wire [63:0] biPassModule_io_dataMem_outputValue_0; // @[AXICache.scala 61:28]
  wire  biPassModule_io_out_valid; // @[AXICache.scala 61:28]
  wire [63:0] biPassModule_io_out_bits_data; // @[AXICache.scala 61:28]
  wire  dataMemory_clock; // @[AXICache.scala 77:26]
  wire  dataMemory_io_read_in_valid; // @[AXICache.scala 77:26]
  wire [31:0] dataMemory_io_read_in_bits_address; // @[AXICache.scala 77:26]
  wire [63:0] dataMemory_io_read_outputValue_0; // @[AXICache.scala 77:26]
  wire  dataMemory_io_write_valid; // @[AXICache.scala 77:26]
  wire [31:0] dataMemory_io_write_bits_address; // @[AXICache.scala 77:26]
  wire [63:0] dataMemory_io_write_bits_inputValue_0; // @[AXICache.scala 77:26]
  wire  metaMemory_clock; // @[AXICache.scala 78:26]
  wire  metaMemory_io_read_in_valid; // @[AXICache.scala 78:26]
  wire  metaMemory_io_read_in_bits_address; // @[AXICache.scala 78:26]
  wire [30:0] metaMemory_io_read_outputValue_0_tag; // @[AXICache.scala 78:26]
  wire [30:0] metaMemory_io_read_outputValue_1_tag; // @[AXICache.scala 78:26]
  wire  metaMemory_io_write_valid; // @[AXICache.scala 78:26]
  wire [1:0] metaMemory_io_write_bits_bank; // @[AXICache.scala 78:26]
  wire  metaMemory_io_write_bits_address; // @[AXICache.scala 78:26]
  wire [30:0] metaMemory_io_write_bits_inputValue_0_tag; // @[AXICache.scala 78:26]
  wire [30:0] metaMemory_io_write_bits_inputValue_1_tag; // @[AXICache.scala 78:26]
  wire  cacheLogic_0_clock; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_reset; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_cpu_req_ready; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_cpu_req_valid; // @[AXICache.scala 81:28]
  wire [31:0] cacheLogic_0_io_cpu_req_bits_addr; // @[AXICache.scala 81:28]
  wire [27:0] cacheLogic_0_io_cpu_req_bits_command; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_0_io_cpu_req_bits_way; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_0_io_cpu_req_bits_replaceWay; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_cpu_resp_valid; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_cpu_resp_bits_iswrite; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_0_io_cpu_resp_bits_way; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_metaMem_write_valid; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_0_io_metaMem_write_bits_bank; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_metaMem_write_bits_address; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_0_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_0_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_validTagBits_write_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_0_io_validTagBits_write_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_validTagBits_write_bits_value; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_validTagBits_read_in_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_0_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_validTagBits_read_out_0; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_validTagBits_read_out_1; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_clock; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_reset; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_io_cpu_req_ready; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_io_cpu_req_valid; // @[AXICache.scala 81:28]
  wire [31:0] cacheLogic_1_io_cpu_req_bits_addr; // @[AXICache.scala 81:28]
  wire [27:0] cacheLogic_1_io_cpu_req_bits_command; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_1_io_cpu_req_bits_way; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_1_io_cpu_req_bits_replaceWay; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_io_cpu_resp_valid; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_io_cpu_resp_bits_iswrite; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_1_io_cpu_resp_bits_way; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_io_metaMem_write_valid; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_1_io_metaMem_write_bits_bank; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_io_metaMem_write_bits_address; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_1_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_1_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_io_validTagBits_write_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_1_io_validTagBits_write_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_io_validTagBits_write_bits_value; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_io_validTagBits_read_in_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_1_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_io_validTagBits_read_out_0; // @[AXICache.scala 81:28]
  wire  cacheLogic_1_io_validTagBits_read_out_1; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_clock; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_reset; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_io_cpu_req_ready; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_io_cpu_req_valid; // @[AXICache.scala 81:28]
  wire [31:0] cacheLogic_2_io_cpu_req_bits_addr; // @[AXICache.scala 81:28]
  wire [27:0] cacheLogic_2_io_cpu_req_bits_command; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_2_io_cpu_req_bits_way; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_2_io_cpu_req_bits_replaceWay; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_io_cpu_resp_valid; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_io_cpu_resp_bits_iswrite; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_2_io_cpu_resp_bits_way; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_io_metaMem_write_valid; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_2_io_metaMem_write_bits_bank; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_io_metaMem_write_bits_address; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_2_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_2_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_io_validTagBits_write_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_2_io_validTagBits_write_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_io_validTagBits_write_bits_value; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_io_validTagBits_read_in_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_2_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_io_validTagBits_read_out_0; // @[AXICache.scala 81:28]
  wire  cacheLogic_2_io_validTagBits_read_out_1; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_clock; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_reset; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_io_cpu_req_ready; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_io_cpu_req_valid; // @[AXICache.scala 81:28]
  wire [31:0] cacheLogic_3_io_cpu_req_bits_addr; // @[AXICache.scala 81:28]
  wire [27:0] cacheLogic_3_io_cpu_req_bits_command; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_3_io_cpu_req_bits_way; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_3_io_cpu_req_bits_replaceWay; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_io_cpu_resp_valid; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_io_cpu_resp_bits_iswrite; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_3_io_cpu_resp_bits_way; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_io_metaMem_write_valid; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_3_io_metaMem_write_bits_bank; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_io_metaMem_write_bits_address; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_3_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_3_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_io_validTagBits_write_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_3_io_validTagBits_write_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_io_validTagBits_write_bits_value; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_io_validTagBits_read_in_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_3_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_io_validTagBits_read_out_0; // @[AXICache.scala 81:28]
  wire  cacheLogic_3_io_validTagBits_read_out_1; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_clock; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_reset; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_io_cpu_req_ready; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_io_cpu_req_valid; // @[AXICache.scala 81:28]
  wire [31:0] cacheLogic_4_io_cpu_req_bits_addr; // @[AXICache.scala 81:28]
  wire [27:0] cacheLogic_4_io_cpu_req_bits_command; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_4_io_cpu_req_bits_way; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_4_io_cpu_req_bits_replaceWay; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_io_cpu_resp_valid; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_io_cpu_resp_bits_iswrite; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_4_io_cpu_resp_bits_way; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_io_metaMem_write_valid; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_4_io_metaMem_write_bits_bank; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_io_metaMem_write_bits_address; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_4_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_4_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_io_validTagBits_write_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_4_io_validTagBits_write_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_io_validTagBits_write_bits_value; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_io_validTagBits_read_in_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_4_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_io_validTagBits_read_out_0; // @[AXICache.scala 81:28]
  wire  cacheLogic_4_io_validTagBits_read_out_1; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_clock; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_reset; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_io_cpu_req_ready; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_io_cpu_req_valid; // @[AXICache.scala 81:28]
  wire [31:0] cacheLogic_5_io_cpu_req_bits_addr; // @[AXICache.scala 81:28]
  wire [27:0] cacheLogic_5_io_cpu_req_bits_command; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_5_io_cpu_req_bits_way; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_5_io_cpu_req_bits_replaceWay; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_io_cpu_resp_valid; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_io_cpu_resp_bits_iswrite; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_5_io_cpu_resp_bits_way; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_io_metaMem_write_valid; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_5_io_metaMem_write_bits_bank; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_io_metaMem_write_bits_address; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_5_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_5_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_io_validTagBits_write_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_5_io_validTagBits_write_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_io_validTagBits_write_bits_value; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_io_validTagBits_read_in_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_5_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_io_validTagBits_read_out_0; // @[AXICache.scala 81:28]
  wire  cacheLogic_5_io_validTagBits_read_out_1; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_clock; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_reset; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_io_cpu_req_ready; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_io_cpu_req_valid; // @[AXICache.scala 81:28]
  wire [31:0] cacheLogic_6_io_cpu_req_bits_addr; // @[AXICache.scala 81:28]
  wire [27:0] cacheLogic_6_io_cpu_req_bits_command; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_6_io_cpu_req_bits_way; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_6_io_cpu_req_bits_replaceWay; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_io_cpu_resp_valid; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_io_cpu_resp_bits_iswrite; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_6_io_cpu_resp_bits_way; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_io_metaMem_write_valid; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_6_io_metaMem_write_bits_bank; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_io_metaMem_write_bits_address; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_6_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_6_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_io_validTagBits_write_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_6_io_validTagBits_write_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_io_validTagBits_write_bits_value; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_io_validTagBits_read_in_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_6_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_io_validTagBits_read_out_0; // @[AXICache.scala 81:28]
  wire  cacheLogic_6_io_validTagBits_read_out_1; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_clock; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_reset; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_io_cpu_req_ready; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_io_cpu_req_valid; // @[AXICache.scala 81:28]
  wire [31:0] cacheLogic_7_io_cpu_req_bits_addr; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_7_io_cpu_req_bits_data; // @[AXICache.scala 81:28]
  wire [27:0] cacheLogic_7_io_cpu_req_bits_command; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_7_io_cpu_req_bits_way; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_7_io_cpu_req_bits_replaceWay; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_io_cpu_resp_valid; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_io_cpu_resp_bits_iswrite; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_7_io_cpu_resp_bits_way; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_io_metaMem_write_valid; // @[AXICache.scala 81:28]
  wire [1:0] cacheLogic_7_io_metaMem_write_bits_bank; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_io_metaMem_write_bits_address; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_7_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 81:28]
  wire [30:0] cacheLogic_7_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_io_dataMem_write_valid; // @[AXICache.scala 81:28]
  wire [31:0] cacheLogic_7_io_dataMem_write_bits_address; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_7_io_dataMem_write_bits_inputValue_0; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_io_validTagBits_write_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_7_io_validTagBits_write_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_io_validTagBits_write_bits_value; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_io_validTagBits_read_in_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_7_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_io_validTagBits_read_out_0; // @[AXICache.scala 81:28]
  wire  cacheLogic_7_io_validTagBits_read_out_1; // @[AXICache.scala 81:28]
  wire  probeUnit_clock; // @[AXICache.scala 85:26]
  wire  probeUnit_reset; // @[AXICache.scala 85:26]
  wire  probeUnit_io_cpu_req_ready; // @[AXICache.scala 85:26]
  wire  probeUnit_io_cpu_req_valid; // @[AXICache.scala 85:26]
  wire [31:0] probeUnit_io_cpu_req_bits_addr; // @[AXICache.scala 85:26]
  wire [27:0] probeUnit_io_cpu_req_bits_command; // @[AXICache.scala 85:26]
  wire  probeUnit_io_cpu_resp_valid; // @[AXICache.scala 85:26]
  wire [1:0] probeUnit_io_cpu_resp_bits_way; // @[AXICache.scala 85:26]
  wire  probeUnit_io_cpu_multiWay_valid; // @[AXICache.scala 85:26]
  wire [1:0] probeUnit_io_cpu_multiWay_bits_way_0; // @[AXICache.scala 85:26]
  wire [1:0] probeUnit_io_cpu_multiWay_bits_way_1; // @[AXICache.scala 85:26]
  wire [31:0] probeUnit_io_cpu_multiWay_bits_addr; // @[AXICache.scala 85:26]
  wire  probeUnit_io_metaMem_read_in_valid; // @[AXICache.scala 85:26]
  wire  probeUnit_io_metaMem_read_in_bits_address; // @[AXICache.scala 85:26]
  wire [30:0] probeUnit_io_metaMem_read_outputValue_0_tag; // @[AXICache.scala 85:26]
  wire [30:0] probeUnit_io_metaMem_read_outputValue_1_tag; // @[AXICache.scala 85:26]
  wire  probeUnit_io_validTagBits_write_valid; // @[AXICache.scala 85:26]
  wire [63:0] probeUnit_io_validTagBits_write_bits_addr; // @[AXICache.scala 85:26]
  wire  probeUnit_io_validTagBits_write_bits_value; // @[AXICache.scala 85:26]
  wire  probeUnit_io_validTagBits_read_in_valid; // @[AXICache.scala 85:26]
  wire [63:0] probeUnit_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 85:26]
  wire  probeUnit_io_validTagBits_read_out_0; // @[AXICache.scala 85:26]
  wire  probeUnit_io_validTagBits_read_out_1; // @[AXICache.scala 85:26]
  wire  validTagBits_clock; // @[AXICache.scala 88:28]
  wire  validTagBits_reset; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_0_write_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_0_write_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_0_write_bits_value; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_0_read_in_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_0_read_in_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_0_read_out_0; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_0_read_out_1; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_1_write_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_1_write_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_1_write_bits_value; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_1_read_in_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_1_read_in_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_1_read_out_0; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_1_read_out_1; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_2_write_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_2_write_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_2_write_bits_value; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_2_read_in_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_2_read_in_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_2_read_out_0; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_2_read_out_1; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_3_write_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_3_write_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_3_write_bits_value; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_3_read_in_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_3_read_in_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_3_read_out_0; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_3_read_out_1; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_4_write_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_4_write_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_4_write_bits_value; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_4_read_in_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_4_read_in_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_4_read_out_0; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_4_read_out_1; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_5_write_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_5_write_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_5_write_bits_value; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_5_read_in_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_5_read_in_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_5_read_out_0; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_5_read_out_1; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_6_write_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_6_write_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_6_write_bits_value; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_6_read_in_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_6_read_in_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_6_read_out_0; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_6_read_out_1; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_7_write_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_7_write_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_7_write_bits_value; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_7_read_in_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_7_read_in_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_7_read_out_0; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_7_read_out_1; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_8_write_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_8_write_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_8_write_bits_value; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_8_read_in_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_8_read_in_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_8_read_out_0; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_8_read_out_1; // @[AXICache.scala 88:28]
  wire  metaWrArb_io_in_0_valid; // @[AXICache.scala 91:27]
  wire [1:0] metaWrArb_io_in_0_bits_bank; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_0_bits_address; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_0_bits_inputValue_0_tag; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_0_bits_inputValue_1_tag; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_1_valid; // @[AXICache.scala 91:27]
  wire [1:0] metaWrArb_io_in_1_bits_bank; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_1_bits_address; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_1_bits_inputValue_0_tag; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_1_bits_inputValue_1_tag; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_2_valid; // @[AXICache.scala 91:27]
  wire [1:0] metaWrArb_io_in_2_bits_bank; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_2_bits_address; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_2_bits_inputValue_0_tag; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_2_bits_inputValue_1_tag; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_3_valid; // @[AXICache.scala 91:27]
  wire [1:0] metaWrArb_io_in_3_bits_bank; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_3_bits_address; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_3_bits_inputValue_0_tag; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_3_bits_inputValue_1_tag; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_4_valid; // @[AXICache.scala 91:27]
  wire [1:0] metaWrArb_io_in_4_bits_bank; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_4_bits_address; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_4_bits_inputValue_0_tag; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_4_bits_inputValue_1_tag; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_5_valid; // @[AXICache.scala 91:27]
  wire [1:0] metaWrArb_io_in_5_bits_bank; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_5_bits_address; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_5_bits_inputValue_0_tag; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_5_bits_inputValue_1_tag; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_6_valid; // @[AXICache.scala 91:27]
  wire [1:0] metaWrArb_io_in_6_bits_bank; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_6_bits_address; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_6_bits_inputValue_0_tag; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_6_bits_inputValue_1_tag; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_7_valid; // @[AXICache.scala 91:27]
  wire [1:0] metaWrArb_io_in_7_bits_bank; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_in_7_bits_address; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_7_bits_inputValue_0_tag; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_in_7_bits_inputValue_1_tag; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_out_valid; // @[AXICache.scala 91:27]
  wire [1:0] metaWrArb_io_out_bits_bank; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_out_bits_address; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_out_bits_inputValue_0_tag; // @[AXICache.scala 91:27]
  wire [30:0] metaWrArb_io_out_bits_inputValue_1_tag; // @[AXICache.scala 91:27]
  bipassLD biPassModule ( // @[AXICache.scala 61:28]
    .clock(biPassModule_clock),
    .reset(biPassModule_reset),
    .io_in_valid(biPassModule_io_in_valid),
    .io_in_bits_addr(biPassModule_io_in_bits_addr),
    .io_in_bits_way(biPassModule_io_in_bits_way),
    .io_dataMem_in_valid(biPassModule_io_dataMem_in_valid),
    .io_dataMem_in_bits_address(biPassModule_io_dataMem_in_bits_address),
    .io_dataMem_outputValue_0(biPassModule_io_dataMem_outputValue_0),
    .io_out_valid(biPassModule_io_out_valid),
    .io_out_bits_data(biPassModule_io_out_bits_data)
  );
  MemBank dataMemory ( // @[AXICache.scala 77:26]
    .clock(dataMemory_clock),
    .io_read_in_valid(dataMemory_io_read_in_valid),
    .io_read_in_bits_address(dataMemory_io_read_in_bits_address),
    .io_read_outputValue_0(dataMemory_io_read_outputValue_0),
    .io_write_valid(dataMemory_io_write_valid),
    .io_write_bits_address(dataMemory_io_write_bits_address),
    .io_write_bits_inputValue_0(dataMemory_io_write_bits_inputValue_0)
  );
  MemBank_1 metaMemory ( // @[AXICache.scala 78:26]
    .clock(metaMemory_clock),
    .io_read_in_valid(metaMemory_io_read_in_valid),
    .io_read_in_bits_address(metaMemory_io_read_in_bits_address),
    .io_read_outputValue_0_tag(metaMemory_io_read_outputValue_0_tag),
    .io_read_outputValue_1_tag(metaMemory_io_read_outputValue_1_tag),
    .io_write_valid(metaMemory_io_write_valid),
    .io_write_bits_bank(metaMemory_io_write_bits_bank),
    .io_write_bits_address(metaMemory_io_write_bits_address),
    .io_write_bits_inputValue_0_tag(metaMemory_io_write_bits_inputValue_0_tag),
    .io_write_bits_inputValue_1_tag(metaMemory_io_write_bits_inputValue_1_tag)
  );
  Gem5CacheLogic cacheLogic_0 ( // @[AXICache.scala 81:28]
    .clock(cacheLogic_0_clock),
    .reset(cacheLogic_0_reset),
    .io_cpu_req_ready(cacheLogic_0_io_cpu_req_ready),
    .io_cpu_req_valid(cacheLogic_0_io_cpu_req_valid),
    .io_cpu_req_bits_addr(cacheLogic_0_io_cpu_req_bits_addr),
    .io_cpu_req_bits_command(cacheLogic_0_io_cpu_req_bits_command),
    .io_cpu_req_bits_way(cacheLogic_0_io_cpu_req_bits_way),
    .io_cpu_req_bits_replaceWay(cacheLogic_0_io_cpu_req_bits_replaceWay),
    .io_cpu_resp_valid(cacheLogic_0_io_cpu_resp_valid),
    .io_cpu_resp_bits_iswrite(cacheLogic_0_io_cpu_resp_bits_iswrite),
    .io_cpu_resp_bits_way(cacheLogic_0_io_cpu_resp_bits_way),
    .io_metaMem_write_valid(cacheLogic_0_io_metaMem_write_valid),
    .io_metaMem_write_bits_bank(cacheLogic_0_io_metaMem_write_bits_bank),
    .io_metaMem_write_bits_address(cacheLogic_0_io_metaMem_write_bits_address),
    .io_metaMem_write_bits_inputValue_0_tag(cacheLogic_0_io_metaMem_write_bits_inputValue_0_tag),
    .io_metaMem_write_bits_inputValue_1_tag(cacheLogic_0_io_metaMem_write_bits_inputValue_1_tag),
    .io_validTagBits_write_valid(cacheLogic_0_io_validTagBits_write_valid),
    .io_validTagBits_write_bits_addr(cacheLogic_0_io_validTagBits_write_bits_addr),
    .io_validTagBits_write_bits_value(cacheLogic_0_io_validTagBits_write_bits_value),
    .io_validTagBits_read_in_valid(cacheLogic_0_io_validTagBits_read_in_valid),
    .io_validTagBits_read_in_bits_addr(cacheLogic_0_io_validTagBits_read_in_bits_addr),
    .io_validTagBits_read_out_0(cacheLogic_0_io_validTagBits_read_out_0),
    .io_validTagBits_read_out_1(cacheLogic_0_io_validTagBits_read_out_1)
  );
  Gem5CacheLogic_1 cacheLogic_1 ( // @[AXICache.scala 81:28]
    .clock(cacheLogic_1_clock),
    .reset(cacheLogic_1_reset),
    .io_cpu_req_ready(cacheLogic_1_io_cpu_req_ready),
    .io_cpu_req_valid(cacheLogic_1_io_cpu_req_valid),
    .io_cpu_req_bits_addr(cacheLogic_1_io_cpu_req_bits_addr),
    .io_cpu_req_bits_command(cacheLogic_1_io_cpu_req_bits_command),
    .io_cpu_req_bits_way(cacheLogic_1_io_cpu_req_bits_way),
    .io_cpu_req_bits_replaceWay(cacheLogic_1_io_cpu_req_bits_replaceWay),
    .io_cpu_resp_valid(cacheLogic_1_io_cpu_resp_valid),
    .io_cpu_resp_bits_iswrite(cacheLogic_1_io_cpu_resp_bits_iswrite),
    .io_cpu_resp_bits_way(cacheLogic_1_io_cpu_resp_bits_way),
    .io_metaMem_write_valid(cacheLogic_1_io_metaMem_write_valid),
    .io_metaMem_write_bits_bank(cacheLogic_1_io_metaMem_write_bits_bank),
    .io_metaMem_write_bits_address(cacheLogic_1_io_metaMem_write_bits_address),
    .io_metaMem_write_bits_inputValue_0_tag(cacheLogic_1_io_metaMem_write_bits_inputValue_0_tag),
    .io_metaMem_write_bits_inputValue_1_tag(cacheLogic_1_io_metaMem_write_bits_inputValue_1_tag),
    .io_validTagBits_write_valid(cacheLogic_1_io_validTagBits_write_valid),
    .io_validTagBits_write_bits_addr(cacheLogic_1_io_validTagBits_write_bits_addr),
    .io_validTagBits_write_bits_value(cacheLogic_1_io_validTagBits_write_bits_value),
    .io_validTagBits_read_in_valid(cacheLogic_1_io_validTagBits_read_in_valid),
    .io_validTagBits_read_in_bits_addr(cacheLogic_1_io_validTagBits_read_in_bits_addr),
    .io_validTagBits_read_out_0(cacheLogic_1_io_validTagBits_read_out_0),
    .io_validTagBits_read_out_1(cacheLogic_1_io_validTagBits_read_out_1)
  );
  Gem5CacheLogic_2 cacheLogic_2 ( // @[AXICache.scala 81:28]
    .clock(cacheLogic_2_clock),
    .reset(cacheLogic_2_reset),
    .io_cpu_req_ready(cacheLogic_2_io_cpu_req_ready),
    .io_cpu_req_valid(cacheLogic_2_io_cpu_req_valid),
    .io_cpu_req_bits_addr(cacheLogic_2_io_cpu_req_bits_addr),
    .io_cpu_req_bits_command(cacheLogic_2_io_cpu_req_bits_command),
    .io_cpu_req_bits_way(cacheLogic_2_io_cpu_req_bits_way),
    .io_cpu_req_bits_replaceWay(cacheLogic_2_io_cpu_req_bits_replaceWay),
    .io_cpu_resp_valid(cacheLogic_2_io_cpu_resp_valid),
    .io_cpu_resp_bits_iswrite(cacheLogic_2_io_cpu_resp_bits_iswrite),
    .io_cpu_resp_bits_way(cacheLogic_2_io_cpu_resp_bits_way),
    .io_metaMem_write_valid(cacheLogic_2_io_metaMem_write_valid),
    .io_metaMem_write_bits_bank(cacheLogic_2_io_metaMem_write_bits_bank),
    .io_metaMem_write_bits_address(cacheLogic_2_io_metaMem_write_bits_address),
    .io_metaMem_write_bits_inputValue_0_tag(cacheLogic_2_io_metaMem_write_bits_inputValue_0_tag),
    .io_metaMem_write_bits_inputValue_1_tag(cacheLogic_2_io_metaMem_write_bits_inputValue_1_tag),
    .io_validTagBits_write_valid(cacheLogic_2_io_validTagBits_write_valid),
    .io_validTagBits_write_bits_addr(cacheLogic_2_io_validTagBits_write_bits_addr),
    .io_validTagBits_write_bits_value(cacheLogic_2_io_validTagBits_write_bits_value),
    .io_validTagBits_read_in_valid(cacheLogic_2_io_validTagBits_read_in_valid),
    .io_validTagBits_read_in_bits_addr(cacheLogic_2_io_validTagBits_read_in_bits_addr),
    .io_validTagBits_read_out_0(cacheLogic_2_io_validTagBits_read_out_0),
    .io_validTagBits_read_out_1(cacheLogic_2_io_validTagBits_read_out_1)
  );
  Gem5CacheLogic_3 cacheLogic_3 ( // @[AXICache.scala 81:28]
    .clock(cacheLogic_3_clock),
    .reset(cacheLogic_3_reset),
    .io_cpu_req_ready(cacheLogic_3_io_cpu_req_ready),
    .io_cpu_req_valid(cacheLogic_3_io_cpu_req_valid),
    .io_cpu_req_bits_addr(cacheLogic_3_io_cpu_req_bits_addr),
    .io_cpu_req_bits_command(cacheLogic_3_io_cpu_req_bits_command),
    .io_cpu_req_bits_way(cacheLogic_3_io_cpu_req_bits_way),
    .io_cpu_req_bits_replaceWay(cacheLogic_3_io_cpu_req_bits_replaceWay),
    .io_cpu_resp_valid(cacheLogic_3_io_cpu_resp_valid),
    .io_cpu_resp_bits_iswrite(cacheLogic_3_io_cpu_resp_bits_iswrite),
    .io_cpu_resp_bits_way(cacheLogic_3_io_cpu_resp_bits_way),
    .io_metaMem_write_valid(cacheLogic_3_io_metaMem_write_valid),
    .io_metaMem_write_bits_bank(cacheLogic_3_io_metaMem_write_bits_bank),
    .io_metaMem_write_bits_address(cacheLogic_3_io_metaMem_write_bits_address),
    .io_metaMem_write_bits_inputValue_0_tag(cacheLogic_3_io_metaMem_write_bits_inputValue_0_tag),
    .io_metaMem_write_bits_inputValue_1_tag(cacheLogic_3_io_metaMem_write_bits_inputValue_1_tag),
    .io_validTagBits_write_valid(cacheLogic_3_io_validTagBits_write_valid),
    .io_validTagBits_write_bits_addr(cacheLogic_3_io_validTagBits_write_bits_addr),
    .io_validTagBits_write_bits_value(cacheLogic_3_io_validTagBits_write_bits_value),
    .io_validTagBits_read_in_valid(cacheLogic_3_io_validTagBits_read_in_valid),
    .io_validTagBits_read_in_bits_addr(cacheLogic_3_io_validTagBits_read_in_bits_addr),
    .io_validTagBits_read_out_0(cacheLogic_3_io_validTagBits_read_out_0),
    .io_validTagBits_read_out_1(cacheLogic_3_io_validTagBits_read_out_1)
  );
  Gem5CacheLogic_4 cacheLogic_4 ( // @[AXICache.scala 81:28]
    .clock(cacheLogic_4_clock),
    .reset(cacheLogic_4_reset),
    .io_cpu_req_ready(cacheLogic_4_io_cpu_req_ready),
    .io_cpu_req_valid(cacheLogic_4_io_cpu_req_valid),
    .io_cpu_req_bits_addr(cacheLogic_4_io_cpu_req_bits_addr),
    .io_cpu_req_bits_command(cacheLogic_4_io_cpu_req_bits_command),
    .io_cpu_req_bits_way(cacheLogic_4_io_cpu_req_bits_way),
    .io_cpu_req_bits_replaceWay(cacheLogic_4_io_cpu_req_bits_replaceWay),
    .io_cpu_resp_valid(cacheLogic_4_io_cpu_resp_valid),
    .io_cpu_resp_bits_iswrite(cacheLogic_4_io_cpu_resp_bits_iswrite),
    .io_cpu_resp_bits_way(cacheLogic_4_io_cpu_resp_bits_way),
    .io_metaMem_write_valid(cacheLogic_4_io_metaMem_write_valid),
    .io_metaMem_write_bits_bank(cacheLogic_4_io_metaMem_write_bits_bank),
    .io_metaMem_write_bits_address(cacheLogic_4_io_metaMem_write_bits_address),
    .io_metaMem_write_bits_inputValue_0_tag(cacheLogic_4_io_metaMem_write_bits_inputValue_0_tag),
    .io_metaMem_write_bits_inputValue_1_tag(cacheLogic_4_io_metaMem_write_bits_inputValue_1_tag),
    .io_validTagBits_write_valid(cacheLogic_4_io_validTagBits_write_valid),
    .io_validTagBits_write_bits_addr(cacheLogic_4_io_validTagBits_write_bits_addr),
    .io_validTagBits_write_bits_value(cacheLogic_4_io_validTagBits_write_bits_value),
    .io_validTagBits_read_in_valid(cacheLogic_4_io_validTagBits_read_in_valid),
    .io_validTagBits_read_in_bits_addr(cacheLogic_4_io_validTagBits_read_in_bits_addr),
    .io_validTagBits_read_out_0(cacheLogic_4_io_validTagBits_read_out_0),
    .io_validTagBits_read_out_1(cacheLogic_4_io_validTagBits_read_out_1)
  );
  Gem5CacheLogic_5 cacheLogic_5 ( // @[AXICache.scala 81:28]
    .clock(cacheLogic_5_clock),
    .reset(cacheLogic_5_reset),
    .io_cpu_req_ready(cacheLogic_5_io_cpu_req_ready),
    .io_cpu_req_valid(cacheLogic_5_io_cpu_req_valid),
    .io_cpu_req_bits_addr(cacheLogic_5_io_cpu_req_bits_addr),
    .io_cpu_req_bits_command(cacheLogic_5_io_cpu_req_bits_command),
    .io_cpu_req_bits_way(cacheLogic_5_io_cpu_req_bits_way),
    .io_cpu_req_bits_replaceWay(cacheLogic_5_io_cpu_req_bits_replaceWay),
    .io_cpu_resp_valid(cacheLogic_5_io_cpu_resp_valid),
    .io_cpu_resp_bits_iswrite(cacheLogic_5_io_cpu_resp_bits_iswrite),
    .io_cpu_resp_bits_way(cacheLogic_5_io_cpu_resp_bits_way),
    .io_metaMem_write_valid(cacheLogic_5_io_metaMem_write_valid),
    .io_metaMem_write_bits_bank(cacheLogic_5_io_metaMem_write_bits_bank),
    .io_metaMem_write_bits_address(cacheLogic_5_io_metaMem_write_bits_address),
    .io_metaMem_write_bits_inputValue_0_tag(cacheLogic_5_io_metaMem_write_bits_inputValue_0_tag),
    .io_metaMem_write_bits_inputValue_1_tag(cacheLogic_5_io_metaMem_write_bits_inputValue_1_tag),
    .io_validTagBits_write_valid(cacheLogic_5_io_validTagBits_write_valid),
    .io_validTagBits_write_bits_addr(cacheLogic_5_io_validTagBits_write_bits_addr),
    .io_validTagBits_write_bits_value(cacheLogic_5_io_validTagBits_write_bits_value),
    .io_validTagBits_read_in_valid(cacheLogic_5_io_validTagBits_read_in_valid),
    .io_validTagBits_read_in_bits_addr(cacheLogic_5_io_validTagBits_read_in_bits_addr),
    .io_validTagBits_read_out_0(cacheLogic_5_io_validTagBits_read_out_0),
    .io_validTagBits_read_out_1(cacheLogic_5_io_validTagBits_read_out_1)
  );
  Gem5CacheLogic_6 cacheLogic_6 ( // @[AXICache.scala 81:28]
    .clock(cacheLogic_6_clock),
    .reset(cacheLogic_6_reset),
    .io_cpu_req_ready(cacheLogic_6_io_cpu_req_ready),
    .io_cpu_req_valid(cacheLogic_6_io_cpu_req_valid),
    .io_cpu_req_bits_addr(cacheLogic_6_io_cpu_req_bits_addr),
    .io_cpu_req_bits_command(cacheLogic_6_io_cpu_req_bits_command),
    .io_cpu_req_bits_way(cacheLogic_6_io_cpu_req_bits_way),
    .io_cpu_req_bits_replaceWay(cacheLogic_6_io_cpu_req_bits_replaceWay),
    .io_cpu_resp_valid(cacheLogic_6_io_cpu_resp_valid),
    .io_cpu_resp_bits_iswrite(cacheLogic_6_io_cpu_resp_bits_iswrite),
    .io_cpu_resp_bits_way(cacheLogic_6_io_cpu_resp_bits_way),
    .io_metaMem_write_valid(cacheLogic_6_io_metaMem_write_valid),
    .io_metaMem_write_bits_bank(cacheLogic_6_io_metaMem_write_bits_bank),
    .io_metaMem_write_bits_address(cacheLogic_6_io_metaMem_write_bits_address),
    .io_metaMem_write_bits_inputValue_0_tag(cacheLogic_6_io_metaMem_write_bits_inputValue_0_tag),
    .io_metaMem_write_bits_inputValue_1_tag(cacheLogic_6_io_metaMem_write_bits_inputValue_1_tag),
    .io_validTagBits_write_valid(cacheLogic_6_io_validTagBits_write_valid),
    .io_validTagBits_write_bits_addr(cacheLogic_6_io_validTagBits_write_bits_addr),
    .io_validTagBits_write_bits_value(cacheLogic_6_io_validTagBits_write_bits_value),
    .io_validTagBits_read_in_valid(cacheLogic_6_io_validTagBits_read_in_valid),
    .io_validTagBits_read_in_bits_addr(cacheLogic_6_io_validTagBits_read_in_bits_addr),
    .io_validTagBits_read_out_0(cacheLogic_6_io_validTagBits_read_out_0),
    .io_validTagBits_read_out_1(cacheLogic_6_io_validTagBits_read_out_1)
  );
  Gem5CacheLogic_7 cacheLogic_7 ( // @[AXICache.scala 81:28]
    .clock(cacheLogic_7_clock),
    .reset(cacheLogic_7_reset),
    .io_cpu_req_ready(cacheLogic_7_io_cpu_req_ready),
    .io_cpu_req_valid(cacheLogic_7_io_cpu_req_valid),
    .io_cpu_req_bits_addr(cacheLogic_7_io_cpu_req_bits_addr),
    .io_cpu_req_bits_data(cacheLogic_7_io_cpu_req_bits_data),
    .io_cpu_req_bits_command(cacheLogic_7_io_cpu_req_bits_command),
    .io_cpu_req_bits_way(cacheLogic_7_io_cpu_req_bits_way),
    .io_cpu_req_bits_replaceWay(cacheLogic_7_io_cpu_req_bits_replaceWay),
    .io_cpu_resp_valid(cacheLogic_7_io_cpu_resp_valid),
    .io_cpu_resp_bits_iswrite(cacheLogic_7_io_cpu_resp_bits_iswrite),
    .io_cpu_resp_bits_way(cacheLogic_7_io_cpu_resp_bits_way),
    .io_metaMem_write_valid(cacheLogic_7_io_metaMem_write_valid),
    .io_metaMem_write_bits_bank(cacheLogic_7_io_metaMem_write_bits_bank),
    .io_metaMem_write_bits_address(cacheLogic_7_io_metaMem_write_bits_address),
    .io_metaMem_write_bits_inputValue_0_tag(cacheLogic_7_io_metaMem_write_bits_inputValue_0_tag),
    .io_metaMem_write_bits_inputValue_1_tag(cacheLogic_7_io_metaMem_write_bits_inputValue_1_tag),
    .io_dataMem_write_valid(cacheLogic_7_io_dataMem_write_valid),
    .io_dataMem_write_bits_address(cacheLogic_7_io_dataMem_write_bits_address),
    .io_dataMem_write_bits_inputValue_0(cacheLogic_7_io_dataMem_write_bits_inputValue_0),
    .io_validTagBits_write_valid(cacheLogic_7_io_validTagBits_write_valid),
    .io_validTagBits_write_bits_addr(cacheLogic_7_io_validTagBits_write_bits_addr),
    .io_validTagBits_write_bits_value(cacheLogic_7_io_validTagBits_write_bits_value),
    .io_validTagBits_read_in_valid(cacheLogic_7_io_validTagBits_read_in_valid),
    .io_validTagBits_read_in_bits_addr(cacheLogic_7_io_validTagBits_read_in_bits_addr),
    .io_validTagBits_read_out_0(cacheLogic_7_io_validTagBits_read_out_0),
    .io_validTagBits_read_out_1(cacheLogic_7_io_validTagBits_read_out_1)
  );
  ProbeUnit probeUnit ( // @[AXICache.scala 85:26]
    .clock(probeUnit_clock),
    .reset(probeUnit_reset),
    .io_cpu_req_ready(probeUnit_io_cpu_req_ready),
    .io_cpu_req_valid(probeUnit_io_cpu_req_valid),
    .io_cpu_req_bits_addr(probeUnit_io_cpu_req_bits_addr),
    .io_cpu_req_bits_command(probeUnit_io_cpu_req_bits_command),
    .io_cpu_resp_valid(probeUnit_io_cpu_resp_valid),
    .io_cpu_resp_bits_way(probeUnit_io_cpu_resp_bits_way),
    .io_cpu_multiWay_valid(probeUnit_io_cpu_multiWay_valid),
    .io_cpu_multiWay_bits_way_0(probeUnit_io_cpu_multiWay_bits_way_0),
    .io_cpu_multiWay_bits_way_1(probeUnit_io_cpu_multiWay_bits_way_1),
    .io_cpu_multiWay_bits_addr(probeUnit_io_cpu_multiWay_bits_addr),
    .io_metaMem_read_in_valid(probeUnit_io_metaMem_read_in_valid),
    .io_metaMem_read_in_bits_address(probeUnit_io_metaMem_read_in_bits_address),
    .io_metaMem_read_outputValue_0_tag(probeUnit_io_metaMem_read_outputValue_0_tag),
    .io_metaMem_read_outputValue_1_tag(probeUnit_io_metaMem_read_outputValue_1_tag),
    .io_validTagBits_write_valid(probeUnit_io_validTagBits_write_valid),
    .io_validTagBits_write_bits_addr(probeUnit_io_validTagBits_write_bits_addr),
    .io_validTagBits_write_bits_value(probeUnit_io_validTagBits_write_bits_value),
    .io_validTagBits_read_in_valid(probeUnit_io_validTagBits_read_in_valid),
    .io_validTagBits_read_in_bits_addr(probeUnit_io_validTagBits_read_in_bits_addr),
    .io_validTagBits_read_out_0(probeUnit_io_validTagBits_read_out_0),
    .io_validTagBits_read_out_1(probeUnit_io_validTagBits_read_out_1)
  );
  paralReg_1 validTagBits ( // @[AXICache.scala 88:28]
    .clock(validTagBits_clock),
    .reset(validTagBits_reset),
    .io_port_0_write_valid(validTagBits_io_port_0_write_valid),
    .io_port_0_write_bits_addr(validTagBits_io_port_0_write_bits_addr),
    .io_port_0_write_bits_value(validTagBits_io_port_0_write_bits_value),
    .io_port_0_read_in_valid(validTagBits_io_port_0_read_in_valid),
    .io_port_0_read_in_bits_addr(validTagBits_io_port_0_read_in_bits_addr),
    .io_port_0_read_out_0(validTagBits_io_port_0_read_out_0),
    .io_port_0_read_out_1(validTagBits_io_port_0_read_out_1),
    .io_port_1_write_valid(validTagBits_io_port_1_write_valid),
    .io_port_1_write_bits_addr(validTagBits_io_port_1_write_bits_addr),
    .io_port_1_write_bits_value(validTagBits_io_port_1_write_bits_value),
    .io_port_1_read_in_valid(validTagBits_io_port_1_read_in_valid),
    .io_port_1_read_in_bits_addr(validTagBits_io_port_1_read_in_bits_addr),
    .io_port_1_read_out_0(validTagBits_io_port_1_read_out_0),
    .io_port_1_read_out_1(validTagBits_io_port_1_read_out_1),
    .io_port_2_write_valid(validTagBits_io_port_2_write_valid),
    .io_port_2_write_bits_addr(validTagBits_io_port_2_write_bits_addr),
    .io_port_2_write_bits_value(validTagBits_io_port_2_write_bits_value),
    .io_port_2_read_in_valid(validTagBits_io_port_2_read_in_valid),
    .io_port_2_read_in_bits_addr(validTagBits_io_port_2_read_in_bits_addr),
    .io_port_2_read_out_0(validTagBits_io_port_2_read_out_0),
    .io_port_2_read_out_1(validTagBits_io_port_2_read_out_1),
    .io_port_3_write_valid(validTagBits_io_port_3_write_valid),
    .io_port_3_write_bits_addr(validTagBits_io_port_3_write_bits_addr),
    .io_port_3_write_bits_value(validTagBits_io_port_3_write_bits_value),
    .io_port_3_read_in_valid(validTagBits_io_port_3_read_in_valid),
    .io_port_3_read_in_bits_addr(validTagBits_io_port_3_read_in_bits_addr),
    .io_port_3_read_out_0(validTagBits_io_port_3_read_out_0),
    .io_port_3_read_out_1(validTagBits_io_port_3_read_out_1),
    .io_port_4_write_valid(validTagBits_io_port_4_write_valid),
    .io_port_4_write_bits_addr(validTagBits_io_port_4_write_bits_addr),
    .io_port_4_write_bits_value(validTagBits_io_port_4_write_bits_value),
    .io_port_4_read_in_valid(validTagBits_io_port_4_read_in_valid),
    .io_port_4_read_in_bits_addr(validTagBits_io_port_4_read_in_bits_addr),
    .io_port_4_read_out_0(validTagBits_io_port_4_read_out_0),
    .io_port_4_read_out_1(validTagBits_io_port_4_read_out_1),
    .io_port_5_write_valid(validTagBits_io_port_5_write_valid),
    .io_port_5_write_bits_addr(validTagBits_io_port_5_write_bits_addr),
    .io_port_5_write_bits_value(validTagBits_io_port_5_write_bits_value),
    .io_port_5_read_in_valid(validTagBits_io_port_5_read_in_valid),
    .io_port_5_read_in_bits_addr(validTagBits_io_port_5_read_in_bits_addr),
    .io_port_5_read_out_0(validTagBits_io_port_5_read_out_0),
    .io_port_5_read_out_1(validTagBits_io_port_5_read_out_1),
    .io_port_6_write_valid(validTagBits_io_port_6_write_valid),
    .io_port_6_write_bits_addr(validTagBits_io_port_6_write_bits_addr),
    .io_port_6_write_bits_value(validTagBits_io_port_6_write_bits_value),
    .io_port_6_read_in_valid(validTagBits_io_port_6_read_in_valid),
    .io_port_6_read_in_bits_addr(validTagBits_io_port_6_read_in_bits_addr),
    .io_port_6_read_out_0(validTagBits_io_port_6_read_out_0),
    .io_port_6_read_out_1(validTagBits_io_port_6_read_out_1),
    .io_port_7_write_valid(validTagBits_io_port_7_write_valid),
    .io_port_7_write_bits_addr(validTagBits_io_port_7_write_bits_addr),
    .io_port_7_write_bits_value(validTagBits_io_port_7_write_bits_value),
    .io_port_7_read_in_valid(validTagBits_io_port_7_read_in_valid),
    .io_port_7_read_in_bits_addr(validTagBits_io_port_7_read_in_bits_addr),
    .io_port_7_read_out_0(validTagBits_io_port_7_read_out_0),
    .io_port_7_read_out_1(validTagBits_io_port_7_read_out_1),
    .io_port_8_write_valid(validTagBits_io_port_8_write_valid),
    .io_port_8_write_bits_addr(validTagBits_io_port_8_write_bits_addr),
    .io_port_8_write_bits_value(validTagBits_io_port_8_write_bits_value),
    .io_port_8_read_in_valid(validTagBits_io_port_8_read_in_valid),
    .io_port_8_read_in_bits_addr(validTagBits_io_port_8_read_in_bits_addr),
    .io_port_8_read_out_0(validTagBits_io_port_8_read_out_0),
    .io_port_8_read_out_1(validTagBits_io_port_8_read_out_1)
  );
  Arbiter_2 metaWrArb ( // @[AXICache.scala 91:27]
    .io_in_0_valid(metaWrArb_io_in_0_valid),
    .io_in_0_bits_bank(metaWrArb_io_in_0_bits_bank),
    .io_in_0_bits_address(metaWrArb_io_in_0_bits_address),
    .io_in_0_bits_inputValue_0_tag(metaWrArb_io_in_0_bits_inputValue_0_tag),
    .io_in_0_bits_inputValue_1_tag(metaWrArb_io_in_0_bits_inputValue_1_tag),
    .io_in_1_valid(metaWrArb_io_in_1_valid),
    .io_in_1_bits_bank(metaWrArb_io_in_1_bits_bank),
    .io_in_1_bits_address(metaWrArb_io_in_1_bits_address),
    .io_in_1_bits_inputValue_0_tag(metaWrArb_io_in_1_bits_inputValue_0_tag),
    .io_in_1_bits_inputValue_1_tag(metaWrArb_io_in_1_bits_inputValue_1_tag),
    .io_in_2_valid(metaWrArb_io_in_2_valid),
    .io_in_2_bits_bank(metaWrArb_io_in_2_bits_bank),
    .io_in_2_bits_address(metaWrArb_io_in_2_bits_address),
    .io_in_2_bits_inputValue_0_tag(metaWrArb_io_in_2_bits_inputValue_0_tag),
    .io_in_2_bits_inputValue_1_tag(metaWrArb_io_in_2_bits_inputValue_1_tag),
    .io_in_3_valid(metaWrArb_io_in_3_valid),
    .io_in_3_bits_bank(metaWrArb_io_in_3_bits_bank),
    .io_in_3_bits_address(metaWrArb_io_in_3_bits_address),
    .io_in_3_bits_inputValue_0_tag(metaWrArb_io_in_3_bits_inputValue_0_tag),
    .io_in_3_bits_inputValue_1_tag(metaWrArb_io_in_3_bits_inputValue_1_tag),
    .io_in_4_valid(metaWrArb_io_in_4_valid),
    .io_in_4_bits_bank(metaWrArb_io_in_4_bits_bank),
    .io_in_4_bits_address(metaWrArb_io_in_4_bits_address),
    .io_in_4_bits_inputValue_0_tag(metaWrArb_io_in_4_bits_inputValue_0_tag),
    .io_in_4_bits_inputValue_1_tag(metaWrArb_io_in_4_bits_inputValue_1_tag),
    .io_in_5_valid(metaWrArb_io_in_5_valid),
    .io_in_5_bits_bank(metaWrArb_io_in_5_bits_bank),
    .io_in_5_bits_address(metaWrArb_io_in_5_bits_address),
    .io_in_5_bits_inputValue_0_tag(metaWrArb_io_in_5_bits_inputValue_0_tag),
    .io_in_5_bits_inputValue_1_tag(metaWrArb_io_in_5_bits_inputValue_1_tag),
    .io_in_6_valid(metaWrArb_io_in_6_valid),
    .io_in_6_bits_bank(metaWrArb_io_in_6_bits_bank),
    .io_in_6_bits_address(metaWrArb_io_in_6_bits_address),
    .io_in_6_bits_inputValue_0_tag(metaWrArb_io_in_6_bits_inputValue_0_tag),
    .io_in_6_bits_inputValue_1_tag(metaWrArb_io_in_6_bits_inputValue_1_tag),
    .io_in_7_valid(metaWrArb_io_in_7_valid),
    .io_in_7_bits_bank(metaWrArb_io_in_7_bits_bank),
    .io_in_7_bits_address(metaWrArb_io_in_7_bits_address),
    .io_in_7_bits_inputValue_0_tag(metaWrArb_io_in_7_bits_inputValue_0_tag),
    .io_in_7_bits_inputValue_1_tag(metaWrArb_io_in_7_bits_inputValue_1_tag),
    .io_out_valid(metaWrArb_io_out_valid),
    .io_out_bits_bank(metaWrArb_io_out_bits_bank),
    .io_out_bits_address(metaWrArb_io_out_bits_address),
    .io_out_bits_inputValue_0_tag(metaWrArb_io_out_bits_inputValue_0_tag),
    .io_out_bits_inputValue_1_tag(metaWrArb_io_out_bits_inputValue_1_tag)
  );
  assign io_cpu_0_resp_valid = cacheLogic_0_io_cpu_resp_valid; // @[AXICache.scala 128:20]
  assign io_cpu_0_resp_bits_iswrite = cacheLogic_0_io_cpu_resp_bits_iswrite; // @[AXICache.scala 128:20]
  assign io_cpu_0_resp_bits_way = cacheLogic_0_io_cpu_resp_bits_way; // @[AXICache.scala 128:20]
  assign io_cpu_1_resp_valid = cacheLogic_1_io_cpu_resp_valid; // @[AXICache.scala 128:20]
  assign io_cpu_1_resp_bits_iswrite = cacheLogic_1_io_cpu_resp_bits_iswrite; // @[AXICache.scala 128:20]
  assign io_cpu_1_resp_bits_way = cacheLogic_1_io_cpu_resp_bits_way; // @[AXICache.scala 128:20]
  assign io_cpu_2_resp_valid = cacheLogic_2_io_cpu_resp_valid; // @[AXICache.scala 128:20]
  assign io_cpu_2_resp_bits_iswrite = cacheLogic_2_io_cpu_resp_bits_iswrite; // @[AXICache.scala 128:20]
  assign io_cpu_2_resp_bits_way = cacheLogic_2_io_cpu_resp_bits_way; // @[AXICache.scala 128:20]
  assign io_cpu_3_resp_valid = cacheLogic_3_io_cpu_resp_valid; // @[AXICache.scala 128:20]
  assign io_cpu_3_resp_bits_iswrite = cacheLogic_3_io_cpu_resp_bits_iswrite; // @[AXICache.scala 128:20]
  assign io_cpu_3_resp_bits_way = cacheLogic_3_io_cpu_resp_bits_way; // @[AXICache.scala 128:20]
  assign io_cpu_4_resp_valid = cacheLogic_4_io_cpu_resp_valid; // @[AXICache.scala 128:20]
  assign io_cpu_4_resp_bits_iswrite = cacheLogic_4_io_cpu_resp_bits_iswrite; // @[AXICache.scala 128:20]
  assign io_cpu_4_resp_bits_way = cacheLogic_4_io_cpu_resp_bits_way; // @[AXICache.scala 128:20]
  assign io_cpu_5_resp_valid = cacheLogic_5_io_cpu_resp_valid; // @[AXICache.scala 128:20]
  assign io_cpu_5_resp_bits_iswrite = cacheLogic_5_io_cpu_resp_bits_iswrite; // @[AXICache.scala 128:20]
  assign io_cpu_5_resp_bits_way = cacheLogic_5_io_cpu_resp_bits_way; // @[AXICache.scala 128:20]
  assign io_cpu_6_resp_valid = cacheLogic_6_io_cpu_resp_valid; // @[AXICache.scala 128:20]
  assign io_cpu_6_resp_bits_iswrite = cacheLogic_6_io_cpu_resp_bits_iswrite; // @[AXICache.scala 128:20]
  assign io_cpu_6_resp_bits_way = cacheLogic_6_io_cpu_resp_bits_way; // @[AXICache.scala 128:20]
  assign io_cpu_7_resp_valid = cacheLogic_7_io_cpu_resp_valid; // @[AXICache.scala 128:20]
  assign io_cpu_7_resp_bits_iswrite = cacheLogic_7_io_cpu_resp_bits_iswrite; // @[AXICache.scala 128:20]
  assign io_cpu_7_resp_bits_way = cacheLogic_7_io_cpu_resp_bits_way; // @[AXICache.scala 128:20]
  assign io_probe_resp_valid = probeUnit_io_cpu_resp_valid; // @[AXICache.scala 133:17]
  assign io_probe_resp_bits_way = probeUnit_io_cpu_resp_bits_way; // @[AXICache.scala 133:17]
  assign io_probe_multiWay_valid = probeUnit_io_cpu_multiWay_valid; // @[AXICache.scala 133:17]
  assign io_probe_multiWay_bits_way_0 = probeUnit_io_cpu_multiWay_bits_way_0; // @[AXICache.scala 133:17]
  assign io_probe_multiWay_bits_way_1 = probeUnit_io_cpu_multiWay_bits_way_1; // @[AXICache.scala 133:17]
  assign io_probe_multiWay_bits_addr = probeUnit_io_cpu_multiWay_bits_addr; // @[AXICache.scala 133:17]
  assign io_bipassLD_out_valid = biPassModule_io_out_valid; // @[AXICache.scala 95:23]
  assign io_bipassLD_out_bits_data = biPassModule_io_out_bits_data; // @[AXICache.scala 95:23]
  assign biPassModule_clock = clock;
  assign biPassModule_reset = reset;
  assign biPassModule_io_in_valid = io_bipassLD_in_valid; // @[AXICache.scala 94:23]
  assign biPassModule_io_in_bits_addr = io_bipassLD_in_bits_addr; // @[AXICache.scala 94:23]
  assign biPassModule_io_in_bits_way = io_bipassLD_in_bits_way; // @[AXICache.scala 94:23]
  assign biPassModule_io_dataMem_outputValue_0 = dataMemory_io_read_outputValue_0; // @[AXICache.scala 97:42]
  assign dataMemory_clock = clock;
  assign dataMemory_io_read_in_valid = biPassModule_io_dataMem_in_valid; // @[AXICache.scala 97:42]
  assign dataMemory_io_read_in_bits_address = biPassModule_io_dataMem_in_bits_address; // @[AXICache.scala 97:42]
  assign dataMemory_io_write_valid = cacheLogic_7_io_dataMem_write_valid; // @[AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35]
  assign dataMemory_io_write_bits_address = cacheLogic_7_io_dataMem_write_bits_address; // @[AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35]
  assign dataMemory_io_write_bits_inputValue_0 = cacheLogic_7_io_dataMem_write_bits_inputValue_0; // @[AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35 AXICache.scala 104:35]
  assign metaMemory_clock = clock;
  assign metaMemory_io_read_in_valid = probeUnit_io_metaMem_read_in_valid; // @[AXICache.scala 98:29]
  assign metaMemory_io_read_in_bits_address = probeUnit_io_metaMem_read_in_bits_address; // @[AXICache.scala 98:29]
  assign metaMemory_io_write_valid = metaWrArb_io_out_valid; // @[AXICache.scala 116:29]
  assign metaMemory_io_write_bits_bank = metaWrArb_io_out_bits_bank; // @[AXICache.scala 113:36]
  assign metaMemory_io_write_bits_address = metaWrArb_io_out_bits_address; // @[AXICache.scala 114:39]
  assign metaMemory_io_write_bits_inputValue_0_tag = metaWrArb_io_out_bits_inputValue_0_tag; // @[AXICache.scala 115:39]
  assign metaMemory_io_write_bits_inputValue_1_tag = metaWrArb_io_out_bits_inputValue_1_tag; // @[AXICache.scala 115:39]
  assign cacheLogic_0_clock = clock;
  assign cacheLogic_0_reset = reset;
  assign cacheLogic_0_io_cpu_req_valid = io_cpu_0_req_valid; // @[AXICache.scala 128:20]
  assign cacheLogic_0_io_cpu_req_bits_addr = io_cpu_0_req_bits_addr; // @[AXICache.scala 128:20]
  assign cacheLogic_0_io_cpu_req_bits_command = io_cpu_0_req_bits_command; // @[AXICache.scala 128:20]
  assign cacheLogic_0_io_cpu_req_bits_way = io_cpu_0_req_bits_way; // @[AXICache.scala 128:20]
  assign cacheLogic_0_io_cpu_req_bits_replaceWay = io_cpu_0_req_bits_replaceWay; // @[AXICache.scala 128:20]
  assign cacheLogic_0_io_validTagBits_read_out_0 = validTagBits_io_port_0_read_out_0; // @[AXICache.scala 127:35]
  assign cacheLogic_0_io_validTagBits_read_out_1 = validTagBits_io_port_0_read_out_1; // @[AXICache.scala 127:35]
  assign cacheLogic_1_clock = clock;
  assign cacheLogic_1_reset = reset;
  assign cacheLogic_1_io_cpu_req_valid = io_cpu_1_req_valid; // @[AXICache.scala 128:20]
  assign cacheLogic_1_io_cpu_req_bits_addr = io_cpu_1_req_bits_addr; // @[AXICache.scala 128:20]
  assign cacheLogic_1_io_cpu_req_bits_command = io_cpu_1_req_bits_command; // @[AXICache.scala 128:20]
  assign cacheLogic_1_io_cpu_req_bits_way = io_cpu_1_req_bits_way; // @[AXICache.scala 128:20]
  assign cacheLogic_1_io_cpu_req_bits_replaceWay = io_cpu_1_req_bits_replaceWay; // @[AXICache.scala 128:20]
  assign cacheLogic_1_io_validTagBits_read_out_0 = validTagBits_io_port_1_read_out_0; // @[AXICache.scala 127:35]
  assign cacheLogic_1_io_validTagBits_read_out_1 = validTagBits_io_port_1_read_out_1; // @[AXICache.scala 127:35]
  assign cacheLogic_2_clock = clock;
  assign cacheLogic_2_reset = reset;
  assign cacheLogic_2_io_cpu_req_valid = io_cpu_2_req_valid; // @[AXICache.scala 128:20]
  assign cacheLogic_2_io_cpu_req_bits_addr = io_cpu_2_req_bits_addr; // @[AXICache.scala 128:20]
  assign cacheLogic_2_io_cpu_req_bits_command = io_cpu_2_req_bits_command; // @[AXICache.scala 128:20]
  assign cacheLogic_2_io_cpu_req_bits_way = io_cpu_2_req_bits_way; // @[AXICache.scala 128:20]
  assign cacheLogic_2_io_cpu_req_bits_replaceWay = io_cpu_2_req_bits_replaceWay; // @[AXICache.scala 128:20]
  assign cacheLogic_2_io_validTagBits_read_out_0 = validTagBits_io_port_2_read_out_0; // @[AXICache.scala 127:35]
  assign cacheLogic_2_io_validTagBits_read_out_1 = validTagBits_io_port_2_read_out_1; // @[AXICache.scala 127:35]
  assign cacheLogic_3_clock = clock;
  assign cacheLogic_3_reset = reset;
  assign cacheLogic_3_io_cpu_req_valid = io_cpu_3_req_valid; // @[AXICache.scala 128:20]
  assign cacheLogic_3_io_cpu_req_bits_addr = io_cpu_3_req_bits_addr; // @[AXICache.scala 128:20]
  assign cacheLogic_3_io_cpu_req_bits_command = io_cpu_3_req_bits_command; // @[AXICache.scala 128:20]
  assign cacheLogic_3_io_cpu_req_bits_way = io_cpu_3_req_bits_way; // @[AXICache.scala 128:20]
  assign cacheLogic_3_io_cpu_req_bits_replaceWay = io_cpu_3_req_bits_replaceWay; // @[AXICache.scala 128:20]
  assign cacheLogic_3_io_validTagBits_read_out_0 = validTagBits_io_port_3_read_out_0; // @[AXICache.scala 127:35]
  assign cacheLogic_3_io_validTagBits_read_out_1 = validTagBits_io_port_3_read_out_1; // @[AXICache.scala 127:35]
  assign cacheLogic_4_clock = clock;
  assign cacheLogic_4_reset = reset;
  assign cacheLogic_4_io_cpu_req_valid = io_cpu_4_req_valid; // @[AXICache.scala 128:20]
  assign cacheLogic_4_io_cpu_req_bits_addr = io_cpu_4_req_bits_addr; // @[AXICache.scala 128:20]
  assign cacheLogic_4_io_cpu_req_bits_command = io_cpu_4_req_bits_command; // @[AXICache.scala 128:20]
  assign cacheLogic_4_io_cpu_req_bits_way = io_cpu_4_req_bits_way; // @[AXICache.scala 128:20]
  assign cacheLogic_4_io_cpu_req_bits_replaceWay = io_cpu_4_req_bits_replaceWay; // @[AXICache.scala 128:20]
  assign cacheLogic_4_io_validTagBits_read_out_0 = validTagBits_io_port_4_read_out_0; // @[AXICache.scala 127:35]
  assign cacheLogic_4_io_validTagBits_read_out_1 = validTagBits_io_port_4_read_out_1; // @[AXICache.scala 127:35]
  assign cacheLogic_5_clock = clock;
  assign cacheLogic_5_reset = reset;
  assign cacheLogic_5_io_cpu_req_valid = io_cpu_5_req_valid; // @[AXICache.scala 128:20]
  assign cacheLogic_5_io_cpu_req_bits_addr = io_cpu_5_req_bits_addr; // @[AXICache.scala 128:20]
  assign cacheLogic_5_io_cpu_req_bits_command = io_cpu_5_req_bits_command; // @[AXICache.scala 128:20]
  assign cacheLogic_5_io_cpu_req_bits_way = io_cpu_5_req_bits_way; // @[AXICache.scala 128:20]
  assign cacheLogic_5_io_cpu_req_bits_replaceWay = io_cpu_5_req_bits_replaceWay; // @[AXICache.scala 128:20]
  assign cacheLogic_5_io_validTagBits_read_out_0 = validTagBits_io_port_5_read_out_0; // @[AXICache.scala 127:35]
  assign cacheLogic_5_io_validTagBits_read_out_1 = validTagBits_io_port_5_read_out_1; // @[AXICache.scala 127:35]
  assign cacheLogic_6_clock = clock;
  assign cacheLogic_6_reset = reset;
  assign cacheLogic_6_io_cpu_req_valid = io_cpu_6_req_valid; // @[AXICache.scala 128:20]
  assign cacheLogic_6_io_cpu_req_bits_addr = io_cpu_6_req_bits_addr; // @[AXICache.scala 128:20]
  assign cacheLogic_6_io_cpu_req_bits_command = io_cpu_6_req_bits_command; // @[AXICache.scala 128:20]
  assign cacheLogic_6_io_cpu_req_bits_way = io_cpu_6_req_bits_way; // @[AXICache.scala 128:20]
  assign cacheLogic_6_io_cpu_req_bits_replaceWay = io_cpu_6_req_bits_replaceWay; // @[AXICache.scala 128:20]
  assign cacheLogic_6_io_validTagBits_read_out_0 = validTagBits_io_port_6_read_out_0; // @[AXICache.scala 127:35]
  assign cacheLogic_6_io_validTagBits_read_out_1 = validTagBits_io_port_6_read_out_1; // @[AXICache.scala 127:35]
  assign cacheLogic_7_clock = clock;
  assign cacheLogic_7_reset = reset;
  assign cacheLogic_7_io_cpu_req_valid = io_cpu_7_req_valid; // @[AXICache.scala 128:20]
  assign cacheLogic_7_io_cpu_req_bits_addr = io_cpu_7_req_bits_addr; // @[AXICache.scala 128:20]
  assign cacheLogic_7_io_cpu_req_bits_data = io_cpu_7_req_bits_data; // @[AXICache.scala 128:20]
  assign cacheLogic_7_io_cpu_req_bits_command = io_cpu_7_req_bits_command; // @[AXICache.scala 128:20]
  assign cacheLogic_7_io_cpu_req_bits_way = io_cpu_7_req_bits_way; // @[AXICache.scala 128:20]
  assign cacheLogic_7_io_cpu_req_bits_replaceWay = io_cpu_7_req_bits_replaceWay; // @[AXICache.scala 128:20]
  assign cacheLogic_7_io_validTagBits_read_out_0 = validTagBits_io_port_7_read_out_0; // @[AXICache.scala 127:35]
  assign cacheLogic_7_io_validTagBits_read_out_1 = validTagBits_io_port_7_read_out_1; // @[AXICache.scala 127:35]
  assign probeUnit_clock = clock;
  assign probeUnit_reset = reset;
  assign probeUnit_io_cpu_req_valid = io_probe_req_valid; // @[AXICache.scala 133:17]
  assign probeUnit_io_cpu_req_bits_addr = io_probe_req_bits_addr; // @[AXICache.scala 133:17]
  assign probeUnit_io_cpu_req_bits_command = io_probe_req_bits_command; // @[AXICache.scala 133:17]
  assign probeUnit_io_metaMem_read_outputValue_0_tag = metaMemory_io_read_outputValue_0_tag; // @[AXICache.scala 98:29]
  assign probeUnit_io_metaMem_read_outputValue_1_tag = metaMemory_io_read_outputValue_1_tag; // @[AXICache.scala 98:29]
  assign probeUnit_io_validTagBits_read_out_0 = validTagBits_io_port_8_read_out_0; // @[AXICache.scala 132:29]
  assign probeUnit_io_validTagBits_read_out_1 = validTagBits_io_port_8_read_out_1; // @[AXICache.scala 132:29]
  assign validTagBits_clock = clock;
  assign validTagBits_reset = reset;
  assign validTagBits_io_port_0_write_valid = cacheLogic_0_io_validTagBits_write_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_0_write_bits_addr = cacheLogic_0_io_validTagBits_write_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_0_write_bits_value = cacheLogic_0_io_validTagBits_write_bits_value; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_0_read_in_valid = cacheLogic_0_io_validTagBits_read_in_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_0_read_in_bits_addr = cacheLogic_0_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_1_write_valid = cacheLogic_1_io_validTagBits_write_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_1_write_bits_addr = cacheLogic_1_io_validTagBits_write_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_1_write_bits_value = cacheLogic_1_io_validTagBits_write_bits_value; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_1_read_in_valid = cacheLogic_1_io_validTagBits_read_in_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_1_read_in_bits_addr = cacheLogic_1_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_2_write_valid = cacheLogic_2_io_validTagBits_write_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_2_write_bits_addr = cacheLogic_2_io_validTagBits_write_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_2_write_bits_value = cacheLogic_2_io_validTagBits_write_bits_value; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_2_read_in_valid = cacheLogic_2_io_validTagBits_read_in_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_2_read_in_bits_addr = cacheLogic_2_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_3_write_valid = cacheLogic_3_io_validTagBits_write_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_3_write_bits_addr = cacheLogic_3_io_validTagBits_write_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_3_write_bits_value = cacheLogic_3_io_validTagBits_write_bits_value; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_3_read_in_valid = cacheLogic_3_io_validTagBits_read_in_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_3_read_in_bits_addr = cacheLogic_3_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_4_write_valid = cacheLogic_4_io_validTagBits_write_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_4_write_bits_addr = cacheLogic_4_io_validTagBits_write_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_4_write_bits_value = cacheLogic_4_io_validTagBits_write_bits_value; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_4_read_in_valid = cacheLogic_4_io_validTagBits_read_in_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_4_read_in_bits_addr = cacheLogic_4_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_5_write_valid = cacheLogic_5_io_validTagBits_write_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_5_write_bits_addr = cacheLogic_5_io_validTagBits_write_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_5_write_bits_value = cacheLogic_5_io_validTagBits_write_bits_value; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_5_read_in_valid = cacheLogic_5_io_validTagBits_read_in_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_5_read_in_bits_addr = cacheLogic_5_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_6_write_valid = cacheLogic_6_io_validTagBits_write_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_6_write_bits_addr = cacheLogic_6_io_validTagBits_write_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_6_write_bits_value = cacheLogic_6_io_validTagBits_write_bits_value; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_6_read_in_valid = cacheLogic_6_io_validTagBits_read_in_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_6_read_in_bits_addr = cacheLogic_6_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_7_write_valid = cacheLogic_7_io_validTagBits_write_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_7_write_bits_addr = cacheLogic_7_io_validTagBits_write_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_7_write_bits_value = cacheLogic_7_io_validTagBits_write_bits_value; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_7_read_in_valid = cacheLogic_7_io_validTagBits_read_in_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_7_read_in_bits_addr = cacheLogic_7_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_8_write_valid = probeUnit_io_validTagBits_write_valid; // @[AXICache.scala 132:29]
  assign validTagBits_io_port_8_write_bits_addr = probeUnit_io_validTagBits_write_bits_addr; // @[AXICache.scala 132:29]
  assign validTagBits_io_port_8_write_bits_value = probeUnit_io_validTagBits_write_bits_value; // @[AXICache.scala 132:29]
  assign validTagBits_io_port_8_read_in_valid = probeUnit_io_validTagBits_read_in_valid; // @[AXICache.scala 132:29]
  assign validTagBits_io_port_8_read_in_bits_addr = probeUnit_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 132:29]
  assign metaWrArb_io_in_0_valid = cacheLogic_0_io_metaMem_write_valid; // @[AXICache.scala 108:33]
  assign metaWrArb_io_in_0_bits_bank = cacheLogic_0_io_metaMem_write_bits_bank; // @[AXICache.scala 105:43]
  assign metaWrArb_io_in_0_bits_address = cacheLogic_0_io_metaMem_write_bits_address; // @[AXICache.scala 106:43]
  assign metaWrArb_io_in_0_bits_inputValue_0_tag = cacheLogic_0_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_0_bits_inputValue_1_tag = cacheLogic_0_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_1_valid = cacheLogic_1_io_metaMem_write_valid; // @[AXICache.scala 108:33]
  assign metaWrArb_io_in_1_bits_bank = cacheLogic_1_io_metaMem_write_bits_bank; // @[AXICache.scala 105:43]
  assign metaWrArb_io_in_1_bits_address = cacheLogic_1_io_metaMem_write_bits_address; // @[AXICache.scala 106:43]
  assign metaWrArb_io_in_1_bits_inputValue_0_tag = cacheLogic_1_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_1_bits_inputValue_1_tag = cacheLogic_1_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_2_valid = cacheLogic_2_io_metaMem_write_valid; // @[AXICache.scala 108:33]
  assign metaWrArb_io_in_2_bits_bank = cacheLogic_2_io_metaMem_write_bits_bank; // @[AXICache.scala 105:43]
  assign metaWrArb_io_in_2_bits_address = cacheLogic_2_io_metaMem_write_bits_address; // @[AXICache.scala 106:43]
  assign metaWrArb_io_in_2_bits_inputValue_0_tag = cacheLogic_2_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_2_bits_inputValue_1_tag = cacheLogic_2_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_3_valid = cacheLogic_3_io_metaMem_write_valid; // @[AXICache.scala 108:33]
  assign metaWrArb_io_in_3_bits_bank = cacheLogic_3_io_metaMem_write_bits_bank; // @[AXICache.scala 105:43]
  assign metaWrArb_io_in_3_bits_address = cacheLogic_3_io_metaMem_write_bits_address; // @[AXICache.scala 106:43]
  assign metaWrArb_io_in_3_bits_inputValue_0_tag = cacheLogic_3_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_3_bits_inputValue_1_tag = cacheLogic_3_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_4_valid = cacheLogic_4_io_metaMem_write_valid; // @[AXICache.scala 108:33]
  assign metaWrArb_io_in_4_bits_bank = cacheLogic_4_io_metaMem_write_bits_bank; // @[AXICache.scala 105:43]
  assign metaWrArb_io_in_4_bits_address = cacheLogic_4_io_metaMem_write_bits_address; // @[AXICache.scala 106:43]
  assign metaWrArb_io_in_4_bits_inputValue_0_tag = cacheLogic_4_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_4_bits_inputValue_1_tag = cacheLogic_4_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_5_valid = cacheLogic_5_io_metaMem_write_valid; // @[AXICache.scala 108:33]
  assign metaWrArb_io_in_5_bits_bank = cacheLogic_5_io_metaMem_write_bits_bank; // @[AXICache.scala 105:43]
  assign metaWrArb_io_in_5_bits_address = cacheLogic_5_io_metaMem_write_bits_address; // @[AXICache.scala 106:43]
  assign metaWrArb_io_in_5_bits_inputValue_0_tag = cacheLogic_5_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_5_bits_inputValue_1_tag = cacheLogic_5_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_6_valid = cacheLogic_6_io_metaMem_write_valid; // @[AXICache.scala 108:33]
  assign metaWrArb_io_in_6_bits_bank = cacheLogic_6_io_metaMem_write_bits_bank; // @[AXICache.scala 105:43]
  assign metaWrArb_io_in_6_bits_address = cacheLogic_6_io_metaMem_write_bits_address; // @[AXICache.scala 106:43]
  assign metaWrArb_io_in_6_bits_inputValue_0_tag = cacheLogic_6_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_6_bits_inputValue_1_tag = cacheLogic_6_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_7_valid = cacheLogic_7_io_metaMem_write_valid; // @[AXICache.scala 108:33]
  assign metaWrArb_io_in_7_bits_bank = cacheLogic_7_io_metaMem_write_bits_bank; // @[AXICache.scala 105:43]
  assign metaWrArb_io_in_7_bits_address = cacheLogic_7_io_metaMem_write_bits_address; // @[AXICache.scala 106:43]
  assign metaWrArb_io_in_7_bits_inputValue_0_tag = cacheLogic_7_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_7_bits_inputValue_1_tag = cacheLogic_7_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 107:43]
endmodule
module FindEmptyLine_9(
  input        io_data_0,
  input        io_data_1,
  input        io_data_2,
  input        io_data_3,
  input        io_data_4,
  input        io_data_5,
  input        io_data_6,
  input        io_data_7,
  input        io_data_8,
  input        io_data_9,
  input        io_data_10,
  input        io_data_11,
  input        io_data_12,
  input        io_data_13,
  input        io_data_14,
  input        io_data_15,
  output [3:0] io_value_bits
);
  wire  _T = ~io_data_0; // @[elements.scala 74:53]
  wire  _T_1 = ~io_data_1; // @[elements.scala 74:53]
  wire  _T_2 = ~io_data_2; // @[elements.scala 74:53]
  wire  _T_3 = ~io_data_3; // @[elements.scala 74:53]
  wire  _T_4 = ~io_data_4; // @[elements.scala 74:53]
  wire  _T_5 = ~io_data_5; // @[elements.scala 74:53]
  wire  _T_6 = ~io_data_6; // @[elements.scala 74:53]
  wire  _T_7 = ~io_data_7; // @[elements.scala 74:53]
  wire  _T_8 = ~io_data_8; // @[elements.scala 74:53]
  wire  _T_9 = ~io_data_9; // @[elements.scala 74:53]
  wire  _T_10 = ~io_data_10; // @[elements.scala 74:53]
  wire  _T_11 = ~io_data_11; // @[elements.scala 74:53]
  wire  _T_12 = ~io_data_12; // @[elements.scala 74:53]
  wire  _T_13 = ~io_data_13; // @[elements.scala 74:53]
  wire  _T_14 = ~io_data_14; // @[elements.scala 74:53]
  wire  _T_15 = ~io_data_15; // @[elements.scala 74:53]
  wire [4:0] _GEN_0 = _T_15 ? 5'hf : 5'h10; // @[elements.scala 74:66]
  wire [4:0] _GEN_2 = _T_14 ? 5'he : _GEN_0; // @[elements.scala 74:66]
  wire [4:0] _GEN_4 = _T_13 ? 5'hd : _GEN_2; // @[elements.scala 74:66]
  wire [4:0] _GEN_6 = _T_12 ? 5'hc : _GEN_4; // @[elements.scala 74:66]
  wire [4:0] _GEN_8 = _T_11 ? 5'hb : _GEN_6; // @[elements.scala 74:66]
  wire [4:0] _GEN_10 = _T_10 ? 5'ha : _GEN_8; // @[elements.scala 74:66]
  wire [4:0] _GEN_12 = _T_9 ? 5'h9 : _GEN_10; // @[elements.scala 74:66]
  wire [4:0] _GEN_14 = _T_8 ? 5'h8 : _GEN_12; // @[elements.scala 74:66]
  wire [4:0] _GEN_16 = _T_7 ? 5'h7 : _GEN_14; // @[elements.scala 74:66]
  wire [4:0] _GEN_18 = _T_6 ? 5'h6 : _GEN_16; // @[elements.scala 74:66]
  wire [4:0] _GEN_20 = _T_5 ? 5'h5 : _GEN_18; // @[elements.scala 74:66]
  wire [4:0] _GEN_22 = _T_4 ? 5'h4 : _GEN_20; // @[elements.scala 74:66]
  wire [4:0] _GEN_24 = _T_3 ? 5'h3 : _GEN_22; // @[elements.scala 74:66]
  wire [4:0] _GEN_26 = _T_2 ? 5'h2 : _GEN_24; // @[elements.scala 74:66]
  wire [4:0] _GEN_28 = _T_1 ? 5'h1 : _GEN_26; // @[elements.scala 74:66]
  wire [4:0] idx = _T ? 5'h0 : _GEN_28; // @[elements.scala 74:66]
  assign io_value_bits = idx[3:0]; // @[elements.scala 79:19]
endmodule
module Find_9(
  input  [31:0] io_key,
  input  [31:0] io_data_0,
  input  [31:0] io_data_1,
  input  [31:0] io_data_2,
  input  [31:0] io_data_3,
  input  [31:0] io_data_4,
  input  [31:0] io_data_5,
  input  [31:0] io_data_6,
  input  [31:0] io_data_7,
  input  [31:0] io_data_8,
  input  [31:0] io_data_9,
  input  [31:0] io_data_10,
  input  [31:0] io_data_11,
  input  [31:0] io_data_12,
  input  [31:0] io_data_13,
  input  [31:0] io_data_14,
  input  [31:0] io_data_15,
  input         io_valid_0,
  input         io_valid_1,
  input         io_valid_2,
  input         io_valid_3,
  input         io_valid_4,
  input         io_valid_5,
  input         io_valid_6,
  input         io_valid_7,
  input         io_valid_8,
  input         io_valid_9,
  input         io_valid_10,
  input         io_valid_11,
  input         io_valid_12,
  input         io_valid_13,
  input         io_valid_14,
  input         io_valid_15,
  output        io_value_valid,
  output [3:0]  io_value_bits
);
  wire  _T = io_data_0 == io_key; // @[elements.scala 35:54]
  wire  _T_1 = io_data_1 == io_key; // @[elements.scala 35:54]
  wire  _T_2 = io_data_2 == io_key; // @[elements.scala 35:54]
  wire  _T_3 = io_data_3 == io_key; // @[elements.scala 35:54]
  wire  _T_4 = io_data_4 == io_key; // @[elements.scala 35:54]
  wire  _T_5 = io_data_5 == io_key; // @[elements.scala 35:54]
  wire  _T_6 = io_data_6 == io_key; // @[elements.scala 35:54]
  wire  _T_7 = io_data_7 == io_key; // @[elements.scala 35:54]
  wire  _T_8 = io_data_8 == io_key; // @[elements.scala 35:54]
  wire  _T_9 = io_data_9 == io_key; // @[elements.scala 35:54]
  wire  _T_10 = io_data_10 == io_key; // @[elements.scala 35:54]
  wire  _T_11 = io_data_11 == io_key; // @[elements.scala 35:54]
  wire  _T_12 = io_data_12 == io_key; // @[elements.scala 35:54]
  wire  _T_13 = io_data_13 == io_key; // @[elements.scala 35:54]
  wire  _T_14 = io_data_14 == io_key; // @[elements.scala 35:54]
  wire  _T_15 = io_data_15 == io_key; // @[elements.scala 35:54]
  wire [7:0] _T_22 = {_T_7,_T_6,_T_5,_T_4,_T_3,_T_2,_T_1,_T}; // @[Cat.scala 29:58]
  wire [15:0] bitmap = {_T_15,_T_14,_T_13,_T_12,_T_11,_T_10,_T_9,_T_8,_T_22}; // @[Cat.scala 29:58]
  wire [7:0] _T_37 = {io_valid_7,io_valid_6,io_valid_5,io_valid_4,io_valid_3,io_valid_2,io_valid_1,io_valid_0}; // @[elements.scala 36:46]
  wire [15:0] _T_45 = {io_valid_15,io_valid_14,io_valid_13,io_valid_12,io_valid_11,io_valid_10,io_valid_9,io_valid_8,_T_37}; // @[elements.scala 36:46]
  wire [15:0] _T_46 = bitmap & _T_45; // @[elements.scala 36:29]
  wire  _T_49 = |_T_46[15:8]; // @[OneHot.scala 32:14]
  wire [7:0] _T_50 = _T_46[15:8] | _T_46[7:0]; // @[OneHot.scala 32:28]
  wire  _T_53 = |_T_50[7:4]; // @[OneHot.scala 32:14]
  wire [3:0] _T_54 = _T_50[7:4] | _T_50[3:0]; // @[OneHot.scala 32:28]
  wire  _T_57 = |_T_54[3:2]; // @[OneHot.scala 32:14]
  wire [1:0] _T_58 = _T_54[3:2] | _T_54[1:0]; // @[OneHot.scala 32:28]
  wire [2:0] _T_61 = {_T_53,_T_57,_T_58[1]}; // @[Cat.scala 29:58]
  assign io_value_valid = _T_46 != 16'h0; // @[elements.scala 39:20]
  assign io_value_bits = {_T_49,_T_61}; // @[elements.scala 38:19]
endmodule
module TBETable(
  input         clock,
  input         reset,
  input         io_write_0_valid,
  input  [63:0] io_write_0_bits_addr,
  input  [1:0]  io_write_0_bits_command,
  input         io_write_0_bits_mask,
  input  [1:0]  io_write_0_bits_inputTBE_state_state,
  input  [2:0]  io_write_0_bits_inputTBE_way,
  input  [31:0] io_write_0_bits_inputTBE_fields_0,
  input         io_write_1_valid,
  input  [63:0] io_write_1_bits_addr,
  input  [1:0]  io_write_1_bits_command,
  input         io_write_1_bits_mask,
  input  [1:0]  io_write_1_bits_inputTBE_state_state,
  input  [2:0]  io_write_1_bits_inputTBE_way,
  input  [31:0] io_write_1_bits_inputTBE_fields_0,
  input         io_write_2_valid,
  input  [63:0] io_write_2_bits_addr,
  input  [1:0]  io_write_2_bits_command,
  input         io_write_2_bits_mask,
  input  [1:0]  io_write_2_bits_inputTBE_state_state,
  input  [2:0]  io_write_2_bits_inputTBE_way,
  input  [31:0] io_write_2_bits_inputTBE_fields_0,
  input         io_write_3_valid,
  input  [63:0] io_write_3_bits_addr,
  input  [1:0]  io_write_3_bits_command,
  input         io_write_3_bits_mask,
  input  [1:0]  io_write_3_bits_inputTBE_state_state,
  input  [2:0]  io_write_3_bits_inputTBE_way,
  input  [31:0] io_write_3_bits_inputTBE_fields_0,
  input         io_write_4_valid,
  input  [63:0] io_write_4_bits_addr,
  input  [1:0]  io_write_4_bits_command,
  input         io_write_4_bits_mask,
  input  [1:0]  io_write_4_bits_inputTBE_state_state,
  input  [2:0]  io_write_4_bits_inputTBE_way,
  input  [31:0] io_write_4_bits_inputTBE_fields_0,
  input         io_write_5_valid,
  input  [63:0] io_write_5_bits_addr,
  input  [1:0]  io_write_5_bits_command,
  input         io_write_5_bits_mask,
  input  [1:0]  io_write_5_bits_inputTBE_state_state,
  input  [2:0]  io_write_5_bits_inputTBE_way,
  input  [31:0] io_write_5_bits_inputTBE_fields_0,
  input         io_write_6_valid,
  input  [63:0] io_write_6_bits_addr,
  input  [1:0]  io_write_6_bits_command,
  input         io_write_6_bits_mask,
  input  [1:0]  io_write_6_bits_inputTBE_state_state,
  input  [2:0]  io_write_6_bits_inputTBE_way,
  input  [31:0] io_write_6_bits_inputTBE_fields_0,
  input         io_write_7_valid,
  input  [63:0] io_write_7_bits_addr,
  input  [1:0]  io_write_7_bits_command,
  input         io_write_7_bits_mask,
  input  [1:0]  io_write_7_bits_inputTBE_state_state,
  input  [2:0]  io_write_7_bits_inputTBE_way,
  input  [31:0] io_write_7_bits_inputTBE_fields_0,
  input         io_read_valid,
  input  [63:0] io_read_bits_addr,
  output [1:0]  io_outputTBE_bits_state_state,
  output [2:0]  io_outputTBE_bits_way,
  output [31:0] io_outputTBE_bits_fields_0,
  output        io_isFull
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
`endif // RANDOMIZE_REG_INIT
  wire  allocLine_io_data_0; // @[TBE.scala 79:25]
  wire  allocLine_io_data_1; // @[TBE.scala 79:25]
  wire  allocLine_io_data_2; // @[TBE.scala 79:25]
  wire  allocLine_io_data_3; // @[TBE.scala 79:25]
  wire  allocLine_io_data_4; // @[TBE.scala 79:25]
  wire  allocLine_io_data_5; // @[TBE.scala 79:25]
  wire  allocLine_io_data_6; // @[TBE.scala 79:25]
  wire  allocLine_io_data_7; // @[TBE.scala 79:25]
  wire  allocLine_io_data_8; // @[TBE.scala 79:25]
  wire  allocLine_io_data_9; // @[TBE.scala 79:25]
  wire  allocLine_io_data_10; // @[TBE.scala 79:25]
  wire  allocLine_io_data_11; // @[TBE.scala 79:25]
  wire  allocLine_io_data_12; // @[TBE.scala 79:25]
  wire  allocLine_io_data_13; // @[TBE.scala 79:25]
  wire  allocLine_io_data_14; // @[TBE.scala 79:25]
  wire  allocLine_io_data_15; // @[TBE.scala 79:25]
  wire [3:0] allocLine_io_value_bits; // @[TBE.scala 79:25]
  wire [31:0] finder_0_io_key; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_0; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_1; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_2; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_3; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_4; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_5; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_6; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_7; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_8; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_9; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_10; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_11; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_12; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_13; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_14; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_15; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_0; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_1; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_2; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_3; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_4; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_5; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_6; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_7; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_8; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_9; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_10; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_11; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_12; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_13; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_14; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_15; // @[TBE.scala 84:24]
  wire  finder_0_io_value_valid; // @[TBE.scala 84:24]
  wire [3:0] finder_0_io_value_bits; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_key; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_0; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_1; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_2; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_3; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_4; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_5; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_6; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_7; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_8; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_9; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_10; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_11; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_12; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_13; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_14; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_15; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_0; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_1; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_2; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_3; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_4; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_5; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_6; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_7; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_8; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_9; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_10; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_11; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_12; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_13; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_14; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_15; // @[TBE.scala 84:24]
  wire  finder_1_io_value_valid; // @[TBE.scala 84:24]
  wire [3:0] finder_1_io_value_bits; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_key; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_0; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_1; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_2; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_3; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_4; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_5; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_6; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_7; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_8; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_9; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_10; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_11; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_12; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_13; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_14; // @[TBE.scala 84:24]
  wire [31:0] finder_2_io_data_15; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_0; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_1; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_2; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_3; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_4; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_5; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_6; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_7; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_8; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_9; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_10; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_11; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_12; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_13; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_14; // @[TBE.scala 84:24]
  wire  finder_2_io_valid_15; // @[TBE.scala 84:24]
  wire  finder_2_io_value_valid; // @[TBE.scala 84:24]
  wire [3:0] finder_2_io_value_bits; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_key; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_0; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_1; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_2; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_3; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_4; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_5; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_6; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_7; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_8; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_9; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_10; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_11; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_12; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_13; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_14; // @[TBE.scala 84:24]
  wire [31:0] finder_3_io_data_15; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_0; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_1; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_2; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_3; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_4; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_5; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_6; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_7; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_8; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_9; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_10; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_11; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_12; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_13; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_14; // @[TBE.scala 84:24]
  wire  finder_3_io_valid_15; // @[TBE.scala 84:24]
  wire  finder_3_io_value_valid; // @[TBE.scala 84:24]
  wire [3:0] finder_3_io_value_bits; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_key; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_0; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_1; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_2; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_3; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_4; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_5; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_6; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_7; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_8; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_9; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_10; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_11; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_12; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_13; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_14; // @[TBE.scala 84:24]
  wire [31:0] finder_4_io_data_15; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_0; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_1; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_2; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_3; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_4; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_5; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_6; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_7; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_8; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_9; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_10; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_11; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_12; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_13; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_14; // @[TBE.scala 84:24]
  wire  finder_4_io_valid_15; // @[TBE.scala 84:24]
  wire  finder_4_io_value_valid; // @[TBE.scala 84:24]
  wire [3:0] finder_4_io_value_bits; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_key; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_0; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_1; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_2; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_3; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_4; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_5; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_6; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_7; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_8; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_9; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_10; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_11; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_12; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_13; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_14; // @[TBE.scala 84:24]
  wire [31:0] finder_5_io_data_15; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_0; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_1; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_2; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_3; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_4; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_5; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_6; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_7; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_8; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_9; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_10; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_11; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_12; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_13; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_14; // @[TBE.scala 84:24]
  wire  finder_5_io_valid_15; // @[TBE.scala 84:24]
  wire  finder_5_io_value_valid; // @[TBE.scala 84:24]
  wire [3:0] finder_5_io_value_bits; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_key; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_0; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_1; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_2; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_3; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_4; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_5; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_6; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_7; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_8; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_9; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_10; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_11; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_12; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_13; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_14; // @[TBE.scala 84:24]
  wire [31:0] finder_6_io_data_15; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_0; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_1; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_2; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_3; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_4; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_5; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_6; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_7; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_8; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_9; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_10; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_11; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_12; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_13; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_14; // @[TBE.scala 84:24]
  wire  finder_6_io_valid_15; // @[TBE.scala 84:24]
  wire  finder_6_io_value_valid; // @[TBE.scala 84:24]
  wire [3:0] finder_6_io_value_bits; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_key; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_0; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_1; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_2; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_3; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_4; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_5; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_6; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_7; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_8; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_9; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_10; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_11; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_12; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_13; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_14; // @[TBE.scala 84:24]
  wire [31:0] finder_7_io_data_15; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_0; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_1; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_2; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_3; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_4; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_5; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_6; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_7; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_8; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_9; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_10; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_11; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_12; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_13; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_14; // @[TBE.scala 84:24]
  wire  finder_7_io_valid_15; // @[TBE.scala 84:24]
  wire  finder_7_io_value_valid; // @[TBE.scala 84:24]
  wire [3:0] finder_7_io_value_bits; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_key; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_0; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_1; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_2; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_3; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_4; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_5; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_6; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_7; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_8; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_9; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_10; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_11; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_12; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_13; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_14; // @[TBE.scala 84:24]
  wire [31:0] finder_8_io_data_15; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_0; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_1; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_2; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_3; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_4; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_5; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_6; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_7; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_8; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_9; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_10; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_11; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_12; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_13; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_14; // @[TBE.scala 84:24]
  wire  finder_8_io_valid_15; // @[TBE.scala 84:24]
  wire  finder_8_io_value_valid; // @[TBE.scala 84:24]
  wire [3:0] finder_8_io_value_bits; // @[TBE.scala 84:24]
  reg [1:0] TBEMemory_0_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_0_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_0_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_1_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_1_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_1_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_2_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_2_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_2_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_3_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_3_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_3_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_4_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_4_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_4_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_5_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_5_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_5_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_6_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_6_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_6_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_7_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_7_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_7_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_8_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_8_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_8_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_9_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_9_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_9_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_10_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_10_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_10_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_11_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_11_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_11_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_12_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_12_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_12_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_13_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_13_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_13_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_14_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_14_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_14_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_15_state_state; // @[TBE.scala 62:26]
  reg [2:0] TBEMemory_15_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_15_fields_0; // @[TBE.scala 62:26]
  reg  TBEValid_0; // @[TBE.scala 63:25]
  reg  TBEValid_1; // @[TBE.scala 63:25]
  reg  TBEValid_2; // @[TBE.scala 63:25]
  reg  TBEValid_3; // @[TBE.scala 63:25]
  reg  TBEValid_4; // @[TBE.scala 63:25]
  reg  TBEValid_5; // @[TBE.scala 63:25]
  reg  TBEValid_6; // @[TBE.scala 63:25]
  reg  TBEValid_7; // @[TBE.scala 63:25]
  reg  TBEValid_8; // @[TBE.scala 63:25]
  reg  TBEValid_9; // @[TBE.scala 63:25]
  reg  TBEValid_10; // @[TBE.scala 63:25]
  reg  TBEValid_11; // @[TBE.scala 63:25]
  reg  TBEValid_12; // @[TBE.scala 63:25]
  reg  TBEValid_13; // @[TBE.scala 63:25]
  reg  TBEValid_14; // @[TBE.scala 63:25]
  reg  TBEValid_15; // @[TBE.scala 63:25]
  reg [31:0] TBEAddr_0; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_1; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_2; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_3; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_4; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_5; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_6; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_7; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_8; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_9; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_10; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_11; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_12; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_13; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_14; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_15; // @[TBE.scala 64:24]
  reg [5:0] counter; // @[TBE.scala 75:24]
  wire [4:0] _T_68 = 5'h10 - 5'h5; // @[TBE.scala 90:40]
  wire [5:0] _GEN_4160 = {{1'd0}, _T_68}; // @[TBE.scala 90:26]
  wire  _T_69 = counter > _GEN_4160; // @[TBE.scala 90:26]
  wire  _T_70 = _T_69 & io_read_valid; // @[TBE.scala 90:58]
  wire  _T_71 = ~finder_8_io_value_valid; // @[TBE.scala 90:69]
  wire  idxReadValid = finder_8_io_value_valid & io_read_valid; // @[TBE.scala 96:50]
  wire [4:0] idxAlloc = {{1'd0}, allocLine_io_value_bits}; // @[TBE.scala 71:22 TBE.scala 81:12]
  wire [31:0] _GEN_0 = 4'h0 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1 = 4'h1 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_1_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2 = 4'h2 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_2_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3 = 4'h3 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_3_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_4 = 4'h4 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_4_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_5 = 4'h5 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_5_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_6 = 4'h6 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_6_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_7 = 4'h7 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_7_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_8 = 4'h8 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_8_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_9 = 4'h9 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_9_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_10 = 4'ha == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_10_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_11 = 4'hb == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_11_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_12 = 4'hc == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_12_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_13 = 4'hd == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_13_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_14 = 4'he == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_14_fields_0; // @[TBE.scala 110:27]
  wire [31:0] _GEN_15 = 4'hf == idxAlloc[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_15_fields_0; // @[TBE.scala 110:27]
  wire [2:0] _GEN_16 = 4'h0 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_0_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_17 = 4'h1 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_1_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_18 = 4'h2 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_2_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_19 = 4'h3 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_3_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_20 = 4'h4 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_4_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_21 = 4'h5 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_5_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_22 = 4'h6 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_6_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_23 = 4'h7 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_7_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_24 = 4'h8 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_8_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_25 = 4'h9 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_9_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_26 = 4'ha == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_10_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_27 = 4'hb == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_11_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_28 = 4'hc == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_12_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_29 = 4'hd == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_13_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_30 = 4'he == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_14_way; // @[TBE.scala 110:27]
  wire [2:0] _GEN_31 = 4'hf == idxAlloc[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_15_way; // @[TBE.scala 110:27]
  wire [1:0] _GEN_32 = 4'h0 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_0_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_33 = 4'h1 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_1_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_34 = 4'h2 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_2_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_35 = 4'h3 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_3_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_36 = 4'h4 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_4_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_37 = 4'h5 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_5_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_38 = 4'h6 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_6_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_39 = 4'h7 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_7_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_40 = 4'h8 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_8_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_41 = 4'h9 == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_9_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_42 = 4'ha == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_10_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_43 = 4'hb == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_11_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_44 = 4'hc == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_12_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_45 = 4'hd == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_13_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_46 = 4'he == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_14_state_state; // @[TBE.scala 110:27]
  wire [1:0] _GEN_47 = 4'hf == idxAlloc[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_15_state_state; // @[TBE.scala 110:27]
  wire [31:0] _GEN_48 = 4'h0 == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_0; // @[TBE.scala 111:25]
  wire [31:0] _GEN_49 = 4'h1 == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_1; // @[TBE.scala 111:25]
  wire [31:0] _GEN_50 = 4'h2 == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_2; // @[TBE.scala 111:25]
  wire [31:0] _GEN_51 = 4'h3 == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_3; // @[TBE.scala 111:25]
  wire [31:0] _GEN_52 = 4'h4 == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_4; // @[TBE.scala 111:25]
  wire [31:0] _GEN_53 = 4'h5 == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_5; // @[TBE.scala 111:25]
  wire [31:0] _GEN_54 = 4'h6 == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_6; // @[TBE.scala 111:25]
  wire [31:0] _GEN_55 = 4'h7 == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_7; // @[TBE.scala 111:25]
  wire [31:0] _GEN_56 = 4'h8 == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_8; // @[TBE.scala 111:25]
  wire [31:0] _GEN_57 = 4'h9 == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_9; // @[TBE.scala 111:25]
  wire [31:0] _GEN_58 = 4'ha == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_10; // @[TBE.scala 111:25]
  wire [31:0] _GEN_59 = 4'hb == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_11; // @[TBE.scala 111:25]
  wire [31:0] _GEN_60 = 4'hc == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_12; // @[TBE.scala 111:25]
  wire [31:0] _GEN_61 = 4'hd == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_13; // @[TBE.scala 111:25]
  wire [31:0] _GEN_62 = 4'he == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_14; // @[TBE.scala 111:25]
  wire [31:0] _GEN_63 = 4'hf == idxAlloc[3:0] ? io_write_0_bits_addr[31:0] : TBEAddr_15; // @[TBE.scala 111:25]
  wire  _GEN_4161 = 4'h0 == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_64 = _GEN_4161 | TBEValid_0; // @[TBE.scala 112:26]
  wire  _GEN_4162 = 4'h1 == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_65 = _GEN_4162 | TBEValid_1; // @[TBE.scala 112:26]
  wire  _GEN_4163 = 4'h2 == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_66 = _GEN_4163 | TBEValid_2; // @[TBE.scala 112:26]
  wire  _GEN_4164 = 4'h3 == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_67 = _GEN_4164 | TBEValid_3; // @[TBE.scala 112:26]
  wire  _GEN_4165 = 4'h4 == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_68 = _GEN_4165 | TBEValid_4; // @[TBE.scala 112:26]
  wire  _GEN_4166 = 4'h5 == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_69 = _GEN_4166 | TBEValid_5; // @[TBE.scala 112:26]
  wire  _GEN_4167 = 4'h6 == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_70 = _GEN_4167 | TBEValid_6; // @[TBE.scala 112:26]
  wire  _GEN_4168 = 4'h7 == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_71 = _GEN_4168 | TBEValid_7; // @[TBE.scala 112:26]
  wire  _GEN_4169 = 4'h8 == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_72 = _GEN_4169 | TBEValid_8; // @[TBE.scala 112:26]
  wire  _GEN_4170 = 4'h9 == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_73 = _GEN_4170 | TBEValid_9; // @[TBE.scala 112:26]
  wire  _GEN_4171 = 4'ha == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_74 = _GEN_4171 | TBEValid_10; // @[TBE.scala 112:26]
  wire  _GEN_4172 = 4'hb == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_75 = _GEN_4172 | TBEValid_11; // @[TBE.scala 112:26]
  wire  _GEN_4173 = 4'hc == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_76 = _GEN_4173 | TBEValid_12; // @[TBE.scala 112:26]
  wire  _GEN_4174 = 4'hd == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_77 = _GEN_4174 | TBEValid_13; // @[TBE.scala 112:26]
  wire  _GEN_4175 = 4'he == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_78 = _GEN_4175 | TBEValid_14; // @[TBE.scala 112:26]
  wire  _GEN_4176 = 4'hf == idxAlloc[3:0]; // @[TBE.scala 112:26]
  wire  _GEN_79 = _GEN_4176 | TBEValid_15; // @[TBE.scala 112:26]
  wire [5:0] _T_88 = counter + 6'h1; // @[TBE.scala 113:26]
  wire  _T_265 = io_write_0_bits_command == 2'h2; // @[TBE.scala 137:46]
  wire  isDealloc_0 = _T_265 & io_write_0_valid; // @[TBE.scala 137:58]
  wire  _T_89 = isDealloc_0 & finder_0_io_value_valid; // @[TBE.scala 114:31]
  wire [4:0] idxUpdate_0 = {{1'd0}, finder_0_io_value_bits}; // @[TBE.scala 73:23 TBE.scala 104:18]
  wire  _GEN_80 = 4'h0 == idxUpdate_0[3:0] ? 1'h0 : TBEValid_0; // @[TBE.scala 115:30]
  wire  _GEN_81 = 4'h1 == idxUpdate_0[3:0] ? 1'h0 : TBEValid_1; // @[TBE.scala 115:30]
  wire  _GEN_82 = 4'h2 == idxUpdate_0[3:0] ? 1'h0 : TBEValid_2; // @[TBE.scala 115:30]
  wire  _GEN_83 = 4'h3 == idxUpdate_0[3:0] ? 1'h0 : TBEValid_3; // @[TBE.scala 115:30]
  wire  _GEN_84 = 4'h4 == idxUpdate_0[3:0] ? 1'h0 : TBEValid_4; // @[TBE.scala 115:30]
  wire  _GEN_85 = 4'h5 == idxUpdate_0[3:0] ? 1'h0 : TBEValid_5; // @[TBE.scala 115:30]
  wire  _GEN_86 = 4'h6 == idxUpdate_0[3:0] ? 1'h0 : TBEValid_6; // @[TBE.scala 115:30]
  wire  _GEN_87 = 4'h7 == idxUpdate_0[3:0] ? 1'h0 : TBEValid_7; // @[TBE.scala 115:30]
  wire  _GEN_88 = 4'h8 == idxUpdate_0[3:0] ? 1'h0 : TBEValid_8; // @[TBE.scala 115:30]
  wire  _GEN_89 = 4'h9 == idxUpdate_0[3:0] ? 1'h0 : TBEValid_9; // @[TBE.scala 115:30]
  wire  _GEN_90 = 4'ha == idxUpdate_0[3:0] ? 1'h0 : TBEValid_10; // @[TBE.scala 115:30]
  wire  _GEN_91 = 4'hb == idxUpdate_0[3:0] ? 1'h0 : TBEValid_11; // @[TBE.scala 115:30]
  wire  _GEN_92 = 4'hc == idxUpdate_0[3:0] ? 1'h0 : TBEValid_12; // @[TBE.scala 115:30]
  wire  _GEN_93 = 4'hd == idxUpdate_0[3:0] ? 1'h0 : TBEValid_13; // @[TBE.scala 115:30]
  wire  _GEN_94 = 4'he == idxUpdate_0[3:0] ? 1'h0 : TBEValid_14; // @[TBE.scala 115:30]
  wire  _GEN_95 = 4'hf == idxUpdate_0[3:0] ? 1'h0 : TBEValid_15; // @[TBE.scala 115:30]
  wire [31:0] _GEN_96 = 4'h0 == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_0_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_97 = 4'h1 == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_1_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_98 = 4'h2 == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_2_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_99 = 4'h3 == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_3_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_100 = 4'h4 == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_4_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_101 = 4'h5 == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_5_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_102 = 4'h6 == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_6_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_103 = 4'h7 == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_7_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_104 = 4'h8 == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_8_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_105 = 4'h9 == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_9_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_106 = 4'ha == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_10_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_107 = 4'hb == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_11_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_108 = 4'hc == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_12_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_109 = 4'hd == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_13_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_110 = 4'he == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_14_fields_0; // @[TBE.scala 116:31]
  wire [31:0] _GEN_111 = 4'hf == idxUpdate_0[3:0] ? 32'h0 : TBEMemory_15_fields_0; // @[TBE.scala 116:31]
  wire [2:0] _GEN_112 = 4'h0 == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_0_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_113 = 4'h1 == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_1_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_114 = 4'h2 == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_2_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_115 = 4'h3 == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_3_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_116 = 4'h4 == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_4_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_117 = 4'h5 == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_5_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_118 = 4'h6 == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_6_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_119 = 4'h7 == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_7_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_120 = 4'h8 == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_8_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_121 = 4'h9 == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_9_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_122 = 4'ha == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_10_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_123 = 4'hb == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_11_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_124 = 4'hc == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_12_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_125 = 4'hd == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_13_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_126 = 4'he == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_14_way; // @[TBE.scala 116:31]
  wire [2:0] _GEN_127 = 4'hf == idxUpdate_0[3:0] ? 3'h2 : TBEMemory_15_way; // @[TBE.scala 116:31]
  wire [1:0] _GEN_128 = 4'h0 == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_0_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_129 = 4'h1 == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_1_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_130 = 4'h2 == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_2_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_131 = 4'h3 == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_3_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_132 = 4'h4 == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_4_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_133 = 4'h5 == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_5_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_134 = 4'h6 == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_6_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_135 = 4'h7 == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_7_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_136 = 4'h8 == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_8_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_137 = 4'h9 == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_9_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_138 = 4'ha == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_10_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_139 = 4'hb == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_11_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_140 = 4'hc == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_12_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_141 = 4'hd == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_13_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_142 = 4'he == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_14_state_state; // @[TBE.scala 116:31]
  wire [1:0] _GEN_143 = 4'hf == idxUpdate_0[3:0] ? 2'h0 : TBEMemory_15_state_state; // @[TBE.scala 116:31]
  wire [31:0] _GEN_144 = 4'h0 == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_0; // @[TBE.scala 117:29]
  wire [31:0] _GEN_145 = 4'h1 == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_1; // @[TBE.scala 117:29]
  wire [31:0] _GEN_146 = 4'h2 == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_2; // @[TBE.scala 117:29]
  wire [31:0] _GEN_147 = 4'h3 == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_3; // @[TBE.scala 117:29]
  wire [31:0] _GEN_148 = 4'h4 == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_4; // @[TBE.scala 117:29]
  wire [31:0] _GEN_149 = 4'h5 == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_5; // @[TBE.scala 117:29]
  wire [31:0] _GEN_150 = 4'h6 == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_6; // @[TBE.scala 117:29]
  wire [31:0] _GEN_151 = 4'h7 == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_7; // @[TBE.scala 117:29]
  wire [31:0] _GEN_152 = 4'h8 == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_8; // @[TBE.scala 117:29]
  wire [31:0] _GEN_153 = 4'h9 == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_9; // @[TBE.scala 117:29]
  wire [31:0] _GEN_154 = 4'ha == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_10; // @[TBE.scala 117:29]
  wire [31:0] _GEN_155 = 4'hb == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_11; // @[TBE.scala 117:29]
  wire [31:0] _GEN_156 = 4'hc == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_12; // @[TBE.scala 117:29]
  wire [31:0] _GEN_157 = 4'hd == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_13; // @[TBE.scala 117:29]
  wire [31:0] _GEN_158 = 4'he == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_14; // @[TBE.scala 117:29]
  wire [31:0] _GEN_159 = 4'hf == idxUpdate_0[3:0] ? 32'h0 : TBEAddr_15; // @[TBE.scala 117:29]
  wire [5:0] _T_96 = counter - 6'h1; // @[TBE.scala 118:26]
  wire  _T_267 = io_write_0_bits_command == 2'h3; // @[TBE.scala 138:44]
  wire  isWrite_0 = _T_267 & io_write_0_valid; // @[TBE.scala 138:55]
  wire  _T_97 = isWrite_0 & finder_0_io_value_valid; // @[TBE.scala 119:29]
  wire  _T_98 = ~io_write_0_bits_mask; // @[TBE.scala 120:35]
  wire [31:0] _GEN_160 = 4'h0 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_161 = 4'h1 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_1_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_162 = 4'h2 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_2_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_163 = 4'h3 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_3_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_164 = 4'h4 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_4_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_165 = 4'h5 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_5_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_166 = 4'h6 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_6_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_167 = 4'h7 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_7_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_168 = 4'h8 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_8_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_169 = 4'h9 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_9_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_170 = 4'ha == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_10_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_171 = 4'hb == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_11_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_172 = 4'hc == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_12_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_173 = 4'hd == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_13_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_174 = 4'he == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_14_fields_0; // @[TBE.scala 121:63]
  wire [31:0] _GEN_175 = 4'hf == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_fields_0 : TBEMemory_15_fields_0; // @[TBE.scala 121:63]
  wire  _T_102 = ~reset; // @[TBE.scala 122:15]
  wire [31:0] _GEN_181 = 4'h1 == idxUpdate_0[3:0] ? TBEMemory_1_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 122:15]
  wire [31:0] _GEN_184 = 4'h2 == idxUpdate_0[3:0] ? TBEMemory_2_fields_0 : _GEN_181; // @[TBE.scala 122:15]
  wire [31:0] _GEN_187 = 4'h3 == idxUpdate_0[3:0] ? TBEMemory_3_fields_0 : _GEN_184; // @[TBE.scala 122:15]
  wire [31:0] _GEN_190 = 4'h4 == idxUpdate_0[3:0] ? TBEMemory_4_fields_0 : _GEN_187; // @[TBE.scala 122:15]
  wire [31:0] _GEN_193 = 4'h5 == idxUpdate_0[3:0] ? TBEMemory_5_fields_0 : _GEN_190; // @[TBE.scala 122:15]
  wire [31:0] _GEN_196 = 4'h6 == idxUpdate_0[3:0] ? TBEMemory_6_fields_0 : _GEN_193; // @[TBE.scala 122:15]
  wire [31:0] _GEN_199 = 4'h7 == idxUpdate_0[3:0] ? TBEMemory_7_fields_0 : _GEN_196; // @[TBE.scala 122:15]
  wire [31:0] _GEN_202 = 4'h8 == idxUpdate_0[3:0] ? TBEMemory_8_fields_0 : _GEN_199; // @[TBE.scala 122:15]
  wire [31:0] _GEN_205 = 4'h9 == idxUpdate_0[3:0] ? TBEMemory_9_fields_0 : _GEN_202; // @[TBE.scala 122:15]
  wire [31:0] _GEN_208 = 4'ha == idxUpdate_0[3:0] ? TBEMemory_10_fields_0 : _GEN_205; // @[TBE.scala 122:15]
  wire [31:0] _GEN_211 = 4'hb == idxUpdate_0[3:0] ? TBEMemory_11_fields_0 : _GEN_208; // @[TBE.scala 122:15]
  wire [31:0] _GEN_214 = 4'hc == idxUpdate_0[3:0] ? TBEMemory_12_fields_0 : _GEN_211; // @[TBE.scala 122:15]
  wire [31:0] _GEN_217 = 4'hd == idxUpdate_0[3:0] ? TBEMemory_13_fields_0 : _GEN_214; // @[TBE.scala 122:15]
  wire [31:0] _GEN_220 = 4'he == idxUpdate_0[3:0] ? TBEMemory_14_fields_0 : _GEN_217; // @[TBE.scala 122:15]
  wire [31:0] _GEN_223 = 4'hf == idxUpdate_0[3:0] ? TBEMemory_15_fields_0 : _GEN_220; // @[TBE.scala 122:15]
  wire [2:0] _GEN_224 = 4'h0 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_0_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_225 = 4'h1 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_1_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_226 = 4'h2 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_2_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_227 = 4'h3 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_3_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_228 = 4'h4 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_4_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_229 = 4'h5 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_5_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_230 = 4'h6 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_6_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_231 = 4'h7 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_7_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_232 = 4'h8 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_8_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_233 = 4'h9 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_9_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_234 = 4'ha == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_10_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_235 = 4'hb == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_11_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_236 = 4'hc == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_12_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_237 = 4'hd == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_13_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_238 = 4'he == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_14_way; // @[TBE.scala 124:37]
  wire [2:0] _GEN_239 = 4'hf == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_way : TBEMemory_15_way; // @[TBE.scala 124:37]
  wire [1:0] _GEN_240 = 4'h0 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_0_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_241 = 4'h1 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_1_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_242 = 4'h2 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_2_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_243 = 4'h3 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_3_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_244 = 4'h4 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_4_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_245 = 4'h5 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_5_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_246 = 4'h6 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_6_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_247 = 4'h7 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_7_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_248 = 4'h8 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_8_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_249 = 4'h9 == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_9_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_250 = 4'ha == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_10_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_251 = 4'hb == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_11_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_252 = 4'hc == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_12_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_253 = 4'hd == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_13_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_254 = 4'he == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_14_state_state; // @[TBE.scala 125:39]
  wire [1:0] _GEN_255 = 4'hf == idxUpdate_0[3:0] ? io_write_0_bits_inputTBE_state_state : TBEMemory_15_state_state; // @[TBE.scala 125:39]
  wire [31:0] _GEN_256 = _T_98 ? _GEN_160 : TBEMemory_0_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_257 = _T_98 ? _GEN_161 : TBEMemory_1_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_258 = _T_98 ? _GEN_162 : TBEMemory_2_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_259 = _T_98 ? _GEN_163 : TBEMemory_3_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_260 = _T_98 ? _GEN_164 : TBEMemory_4_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_261 = _T_98 ? _GEN_165 : TBEMemory_5_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_262 = _T_98 ? _GEN_166 : TBEMemory_6_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_263 = _T_98 ? _GEN_167 : TBEMemory_7_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_264 = _T_98 ? _GEN_168 : TBEMemory_8_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_265 = _T_98 ? _GEN_169 : TBEMemory_9_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_266 = _T_98 ? _GEN_170 : TBEMemory_10_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_267 = _T_98 ? _GEN_171 : TBEMemory_11_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_268 = _T_98 ? _GEN_172 : TBEMemory_12_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_269 = _T_98 ? _GEN_173 : TBEMemory_13_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_270 = _T_98 ? _GEN_174 : TBEMemory_14_fields_0; // @[TBE.scala 120:53]
  wire [31:0] _GEN_271 = _T_98 ? _GEN_175 : TBEMemory_15_fields_0; // @[TBE.scala 120:53]
  wire [2:0] _GEN_272 = _T_98 ? TBEMemory_0_way : _GEN_224; // @[TBE.scala 120:53]
  wire [2:0] _GEN_273 = _T_98 ? TBEMemory_1_way : _GEN_225; // @[TBE.scala 120:53]
  wire [2:0] _GEN_274 = _T_98 ? TBEMemory_2_way : _GEN_226; // @[TBE.scala 120:53]
  wire [2:0] _GEN_275 = _T_98 ? TBEMemory_3_way : _GEN_227; // @[TBE.scala 120:53]
  wire [2:0] _GEN_276 = _T_98 ? TBEMemory_4_way : _GEN_228; // @[TBE.scala 120:53]
  wire [2:0] _GEN_277 = _T_98 ? TBEMemory_5_way : _GEN_229; // @[TBE.scala 120:53]
  wire [2:0] _GEN_278 = _T_98 ? TBEMemory_6_way : _GEN_230; // @[TBE.scala 120:53]
  wire [2:0] _GEN_279 = _T_98 ? TBEMemory_7_way : _GEN_231; // @[TBE.scala 120:53]
  wire [2:0] _GEN_280 = _T_98 ? TBEMemory_8_way : _GEN_232; // @[TBE.scala 120:53]
  wire [2:0] _GEN_281 = _T_98 ? TBEMemory_9_way : _GEN_233; // @[TBE.scala 120:53]
  wire [2:0] _GEN_282 = _T_98 ? TBEMemory_10_way : _GEN_234; // @[TBE.scala 120:53]
  wire [2:0] _GEN_283 = _T_98 ? TBEMemory_11_way : _GEN_235; // @[TBE.scala 120:53]
  wire [2:0] _GEN_284 = _T_98 ? TBEMemory_12_way : _GEN_236; // @[TBE.scala 120:53]
  wire [2:0] _GEN_285 = _T_98 ? TBEMemory_13_way : _GEN_237; // @[TBE.scala 120:53]
  wire [2:0] _GEN_286 = _T_98 ? TBEMemory_14_way : _GEN_238; // @[TBE.scala 120:53]
  wire [2:0] _GEN_287 = _T_98 ? TBEMemory_15_way : _GEN_239; // @[TBE.scala 120:53]
  wire [1:0] _GEN_288 = _T_98 ? TBEMemory_0_state_state : _GEN_240; // @[TBE.scala 120:53]
  wire [1:0] _GEN_289 = _T_98 ? TBEMemory_1_state_state : _GEN_241; // @[TBE.scala 120:53]
  wire [1:0] _GEN_290 = _T_98 ? TBEMemory_2_state_state : _GEN_242; // @[TBE.scala 120:53]
  wire [1:0] _GEN_291 = _T_98 ? TBEMemory_3_state_state : _GEN_243; // @[TBE.scala 120:53]
  wire [1:0] _GEN_292 = _T_98 ? TBEMemory_4_state_state : _GEN_244; // @[TBE.scala 120:53]
  wire [1:0] _GEN_293 = _T_98 ? TBEMemory_5_state_state : _GEN_245; // @[TBE.scala 120:53]
  wire [1:0] _GEN_294 = _T_98 ? TBEMemory_6_state_state : _GEN_246; // @[TBE.scala 120:53]
  wire [1:0] _GEN_295 = _T_98 ? TBEMemory_7_state_state : _GEN_247; // @[TBE.scala 120:53]
  wire [1:0] _GEN_296 = _T_98 ? TBEMemory_8_state_state : _GEN_248; // @[TBE.scala 120:53]
  wire [1:0] _GEN_297 = _T_98 ? TBEMemory_9_state_state : _GEN_249; // @[TBE.scala 120:53]
  wire [1:0] _GEN_298 = _T_98 ? TBEMemory_10_state_state : _GEN_250; // @[TBE.scala 120:53]
  wire [1:0] _GEN_299 = _T_98 ? TBEMemory_11_state_state : _GEN_251; // @[TBE.scala 120:53]
  wire [1:0] _GEN_300 = _T_98 ? TBEMemory_12_state_state : _GEN_252; // @[TBE.scala 120:53]
  wire [1:0] _GEN_301 = _T_98 ? TBEMemory_13_state_state : _GEN_253; // @[TBE.scala 120:53]
  wire [1:0] _GEN_302 = _T_98 ? TBEMemory_14_state_state : _GEN_254; // @[TBE.scala 120:53]
  wire [1:0] _GEN_303 = _T_98 ? TBEMemory_15_state_state : _GEN_255; // @[TBE.scala 120:53]
  wire [31:0] _GEN_304 = _T_97 ? _GEN_256 : TBEMemory_0_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_305 = _T_97 ? _GEN_257 : TBEMemory_1_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_306 = _T_97 ? _GEN_258 : TBEMemory_2_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_307 = _T_97 ? _GEN_259 : TBEMemory_3_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_308 = _T_97 ? _GEN_260 : TBEMemory_4_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_309 = _T_97 ? _GEN_261 : TBEMemory_5_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_310 = _T_97 ? _GEN_262 : TBEMemory_6_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_311 = _T_97 ? _GEN_263 : TBEMemory_7_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_312 = _T_97 ? _GEN_264 : TBEMemory_8_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_313 = _T_97 ? _GEN_265 : TBEMemory_9_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_314 = _T_97 ? _GEN_266 : TBEMemory_10_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_315 = _T_97 ? _GEN_267 : TBEMemory_11_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_316 = _T_97 ? _GEN_268 : TBEMemory_12_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_317 = _T_97 ? _GEN_269 : TBEMemory_13_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_318 = _T_97 ? _GEN_270 : TBEMemory_14_fields_0; // @[TBE.scala 119:57]
  wire [31:0] _GEN_319 = _T_97 ? _GEN_271 : TBEMemory_15_fields_0; // @[TBE.scala 119:57]
  wire [2:0] _GEN_320 = _T_97 ? _GEN_272 : TBEMemory_0_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_321 = _T_97 ? _GEN_273 : TBEMemory_1_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_322 = _T_97 ? _GEN_274 : TBEMemory_2_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_323 = _T_97 ? _GEN_275 : TBEMemory_3_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_324 = _T_97 ? _GEN_276 : TBEMemory_4_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_325 = _T_97 ? _GEN_277 : TBEMemory_5_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_326 = _T_97 ? _GEN_278 : TBEMemory_6_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_327 = _T_97 ? _GEN_279 : TBEMemory_7_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_328 = _T_97 ? _GEN_280 : TBEMemory_8_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_329 = _T_97 ? _GEN_281 : TBEMemory_9_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_330 = _T_97 ? _GEN_282 : TBEMemory_10_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_331 = _T_97 ? _GEN_283 : TBEMemory_11_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_332 = _T_97 ? _GEN_284 : TBEMemory_12_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_333 = _T_97 ? _GEN_285 : TBEMemory_13_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_334 = _T_97 ? _GEN_286 : TBEMemory_14_way; // @[TBE.scala 119:57]
  wire [2:0] _GEN_335 = _T_97 ? _GEN_287 : TBEMemory_15_way; // @[TBE.scala 119:57]
  wire [1:0] _GEN_336 = _T_97 ? _GEN_288 : TBEMemory_0_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_337 = _T_97 ? _GEN_289 : TBEMemory_1_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_338 = _T_97 ? _GEN_290 : TBEMemory_2_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_339 = _T_97 ? _GEN_291 : TBEMemory_3_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_340 = _T_97 ? _GEN_292 : TBEMemory_4_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_341 = _T_97 ? _GEN_293 : TBEMemory_5_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_342 = _T_97 ? _GEN_294 : TBEMemory_6_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_343 = _T_97 ? _GEN_295 : TBEMemory_7_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_344 = _T_97 ? _GEN_296 : TBEMemory_8_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_345 = _T_97 ? _GEN_297 : TBEMemory_9_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_346 = _T_97 ? _GEN_298 : TBEMemory_10_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_347 = _T_97 ? _GEN_299 : TBEMemory_11_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_348 = _T_97 ? _GEN_300 : TBEMemory_12_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_349 = _T_97 ? _GEN_301 : TBEMemory_13_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_350 = _T_97 ? _GEN_302 : TBEMemory_14_state_state; // @[TBE.scala 119:57]
  wire [1:0] _GEN_351 = _T_97 ? _GEN_303 : TBEMemory_15_state_state; // @[TBE.scala 119:57]
  wire  _GEN_352 = _T_89 ? _GEN_80 : TBEValid_0; // @[TBE.scala 114:59]
  wire  _GEN_353 = _T_89 ? _GEN_81 : TBEValid_1; // @[TBE.scala 114:59]
  wire  _GEN_354 = _T_89 ? _GEN_82 : TBEValid_2; // @[TBE.scala 114:59]
  wire  _GEN_355 = _T_89 ? _GEN_83 : TBEValid_3; // @[TBE.scala 114:59]
  wire  _GEN_356 = _T_89 ? _GEN_84 : TBEValid_4; // @[TBE.scala 114:59]
  wire  _GEN_357 = _T_89 ? _GEN_85 : TBEValid_5; // @[TBE.scala 114:59]
  wire  _GEN_358 = _T_89 ? _GEN_86 : TBEValid_6; // @[TBE.scala 114:59]
  wire  _GEN_359 = _T_89 ? _GEN_87 : TBEValid_7; // @[TBE.scala 114:59]
  wire  _GEN_360 = _T_89 ? _GEN_88 : TBEValid_8; // @[TBE.scala 114:59]
  wire  _GEN_361 = _T_89 ? _GEN_89 : TBEValid_9; // @[TBE.scala 114:59]
  wire  _GEN_362 = _T_89 ? _GEN_90 : TBEValid_10; // @[TBE.scala 114:59]
  wire  _GEN_363 = _T_89 ? _GEN_91 : TBEValid_11; // @[TBE.scala 114:59]
  wire  _GEN_364 = _T_89 ? _GEN_92 : TBEValid_12; // @[TBE.scala 114:59]
  wire  _GEN_365 = _T_89 ? _GEN_93 : TBEValid_13; // @[TBE.scala 114:59]
  wire  _GEN_366 = _T_89 ? _GEN_94 : TBEValid_14; // @[TBE.scala 114:59]
  wire  _GEN_367 = _T_89 ? _GEN_95 : TBEValid_15; // @[TBE.scala 114:59]
  wire [31:0] _GEN_368 = _T_89 ? _GEN_96 : _GEN_304; // @[TBE.scala 114:59]
  wire [31:0] _GEN_369 = _T_89 ? _GEN_97 : _GEN_305; // @[TBE.scala 114:59]
  wire [31:0] _GEN_370 = _T_89 ? _GEN_98 : _GEN_306; // @[TBE.scala 114:59]
  wire [31:0] _GEN_371 = _T_89 ? _GEN_99 : _GEN_307; // @[TBE.scala 114:59]
  wire [31:0] _GEN_372 = _T_89 ? _GEN_100 : _GEN_308; // @[TBE.scala 114:59]
  wire [31:0] _GEN_373 = _T_89 ? _GEN_101 : _GEN_309; // @[TBE.scala 114:59]
  wire [31:0] _GEN_374 = _T_89 ? _GEN_102 : _GEN_310; // @[TBE.scala 114:59]
  wire [31:0] _GEN_375 = _T_89 ? _GEN_103 : _GEN_311; // @[TBE.scala 114:59]
  wire [31:0] _GEN_376 = _T_89 ? _GEN_104 : _GEN_312; // @[TBE.scala 114:59]
  wire [31:0] _GEN_377 = _T_89 ? _GEN_105 : _GEN_313; // @[TBE.scala 114:59]
  wire [31:0] _GEN_378 = _T_89 ? _GEN_106 : _GEN_314; // @[TBE.scala 114:59]
  wire [31:0] _GEN_379 = _T_89 ? _GEN_107 : _GEN_315; // @[TBE.scala 114:59]
  wire [31:0] _GEN_380 = _T_89 ? _GEN_108 : _GEN_316; // @[TBE.scala 114:59]
  wire [31:0] _GEN_381 = _T_89 ? _GEN_109 : _GEN_317; // @[TBE.scala 114:59]
  wire [31:0] _GEN_382 = _T_89 ? _GEN_110 : _GEN_318; // @[TBE.scala 114:59]
  wire [31:0] _GEN_383 = _T_89 ? _GEN_111 : _GEN_319; // @[TBE.scala 114:59]
  wire [2:0] _GEN_384 = _T_89 ? _GEN_112 : _GEN_320; // @[TBE.scala 114:59]
  wire [2:0] _GEN_385 = _T_89 ? _GEN_113 : _GEN_321; // @[TBE.scala 114:59]
  wire [2:0] _GEN_386 = _T_89 ? _GEN_114 : _GEN_322; // @[TBE.scala 114:59]
  wire [2:0] _GEN_387 = _T_89 ? _GEN_115 : _GEN_323; // @[TBE.scala 114:59]
  wire [2:0] _GEN_388 = _T_89 ? _GEN_116 : _GEN_324; // @[TBE.scala 114:59]
  wire [2:0] _GEN_389 = _T_89 ? _GEN_117 : _GEN_325; // @[TBE.scala 114:59]
  wire [2:0] _GEN_390 = _T_89 ? _GEN_118 : _GEN_326; // @[TBE.scala 114:59]
  wire [2:0] _GEN_391 = _T_89 ? _GEN_119 : _GEN_327; // @[TBE.scala 114:59]
  wire [2:0] _GEN_392 = _T_89 ? _GEN_120 : _GEN_328; // @[TBE.scala 114:59]
  wire [2:0] _GEN_393 = _T_89 ? _GEN_121 : _GEN_329; // @[TBE.scala 114:59]
  wire [2:0] _GEN_394 = _T_89 ? _GEN_122 : _GEN_330; // @[TBE.scala 114:59]
  wire [2:0] _GEN_395 = _T_89 ? _GEN_123 : _GEN_331; // @[TBE.scala 114:59]
  wire [2:0] _GEN_396 = _T_89 ? _GEN_124 : _GEN_332; // @[TBE.scala 114:59]
  wire [2:0] _GEN_397 = _T_89 ? _GEN_125 : _GEN_333; // @[TBE.scala 114:59]
  wire [2:0] _GEN_398 = _T_89 ? _GEN_126 : _GEN_334; // @[TBE.scala 114:59]
  wire [2:0] _GEN_399 = _T_89 ? _GEN_127 : _GEN_335; // @[TBE.scala 114:59]
  wire [1:0] _GEN_400 = _T_89 ? _GEN_128 : _GEN_336; // @[TBE.scala 114:59]
  wire [1:0] _GEN_401 = _T_89 ? _GEN_129 : _GEN_337; // @[TBE.scala 114:59]
  wire [1:0] _GEN_402 = _T_89 ? _GEN_130 : _GEN_338; // @[TBE.scala 114:59]
  wire [1:0] _GEN_403 = _T_89 ? _GEN_131 : _GEN_339; // @[TBE.scala 114:59]
  wire [1:0] _GEN_404 = _T_89 ? _GEN_132 : _GEN_340; // @[TBE.scala 114:59]
  wire [1:0] _GEN_405 = _T_89 ? _GEN_133 : _GEN_341; // @[TBE.scala 114:59]
  wire [1:0] _GEN_406 = _T_89 ? _GEN_134 : _GEN_342; // @[TBE.scala 114:59]
  wire [1:0] _GEN_407 = _T_89 ? _GEN_135 : _GEN_343; // @[TBE.scala 114:59]
  wire [1:0] _GEN_408 = _T_89 ? _GEN_136 : _GEN_344; // @[TBE.scala 114:59]
  wire [1:0] _GEN_409 = _T_89 ? _GEN_137 : _GEN_345; // @[TBE.scala 114:59]
  wire [1:0] _GEN_410 = _T_89 ? _GEN_138 : _GEN_346; // @[TBE.scala 114:59]
  wire [1:0] _GEN_411 = _T_89 ? _GEN_139 : _GEN_347; // @[TBE.scala 114:59]
  wire [1:0] _GEN_412 = _T_89 ? _GEN_140 : _GEN_348; // @[TBE.scala 114:59]
  wire [1:0] _GEN_413 = _T_89 ? _GEN_141 : _GEN_349; // @[TBE.scala 114:59]
  wire [1:0] _GEN_414 = _T_89 ? _GEN_142 : _GEN_350; // @[TBE.scala 114:59]
  wire [1:0] _GEN_415 = _T_89 ? _GEN_143 : _GEN_351; // @[TBE.scala 114:59]
  wire [31:0] _GEN_416 = _T_89 ? _GEN_144 : TBEAddr_0; // @[TBE.scala 114:59]
  wire [31:0] _GEN_417 = _T_89 ? _GEN_145 : TBEAddr_1; // @[TBE.scala 114:59]
  wire [31:0] _GEN_418 = _T_89 ? _GEN_146 : TBEAddr_2; // @[TBE.scala 114:59]
  wire [31:0] _GEN_419 = _T_89 ? _GEN_147 : TBEAddr_3; // @[TBE.scala 114:59]
  wire [31:0] _GEN_420 = _T_89 ? _GEN_148 : TBEAddr_4; // @[TBE.scala 114:59]
  wire [31:0] _GEN_421 = _T_89 ? _GEN_149 : TBEAddr_5; // @[TBE.scala 114:59]
  wire [31:0] _GEN_422 = _T_89 ? _GEN_150 : TBEAddr_6; // @[TBE.scala 114:59]
  wire [31:0] _GEN_423 = _T_89 ? _GEN_151 : TBEAddr_7; // @[TBE.scala 114:59]
  wire [31:0] _GEN_424 = _T_89 ? _GEN_152 : TBEAddr_8; // @[TBE.scala 114:59]
  wire [31:0] _GEN_425 = _T_89 ? _GEN_153 : TBEAddr_9; // @[TBE.scala 114:59]
  wire [31:0] _GEN_426 = _T_89 ? _GEN_154 : TBEAddr_10; // @[TBE.scala 114:59]
  wire [31:0] _GEN_427 = _T_89 ? _GEN_155 : TBEAddr_11; // @[TBE.scala 114:59]
  wire [31:0] _GEN_428 = _T_89 ? _GEN_156 : TBEAddr_12; // @[TBE.scala 114:59]
  wire [31:0] _GEN_429 = _T_89 ? _GEN_157 : TBEAddr_13; // @[TBE.scala 114:59]
  wire [31:0] _GEN_430 = _T_89 ? _GEN_158 : TBEAddr_14; // @[TBE.scala 114:59]
  wire [31:0] _GEN_431 = _T_89 ? _GEN_159 : TBEAddr_15; // @[TBE.scala 114:59]
  wire  _T_263 = io_write_0_bits_command == 2'h1; // @[TBE.scala 136:44]
  wire  isAlloc_0 = _T_263 & io_write_0_valid; // @[TBE.scala 136:54]
  wire [31:0] _GEN_433 = isAlloc_0 ? _GEN_0 : _GEN_368; // @[TBE.scala 109:24]
  wire [31:0] _GEN_434 = isAlloc_0 ? _GEN_1 : _GEN_369; // @[TBE.scala 109:24]
  wire [31:0] _GEN_435 = isAlloc_0 ? _GEN_2 : _GEN_370; // @[TBE.scala 109:24]
  wire [31:0] _GEN_436 = isAlloc_0 ? _GEN_3 : _GEN_371; // @[TBE.scala 109:24]
  wire [31:0] _GEN_437 = isAlloc_0 ? _GEN_4 : _GEN_372; // @[TBE.scala 109:24]
  wire [31:0] _GEN_438 = isAlloc_0 ? _GEN_5 : _GEN_373; // @[TBE.scala 109:24]
  wire [31:0] _GEN_439 = isAlloc_0 ? _GEN_6 : _GEN_374; // @[TBE.scala 109:24]
  wire [31:0] _GEN_440 = isAlloc_0 ? _GEN_7 : _GEN_375; // @[TBE.scala 109:24]
  wire [31:0] _GEN_441 = isAlloc_0 ? _GEN_8 : _GEN_376; // @[TBE.scala 109:24]
  wire [31:0] _GEN_442 = isAlloc_0 ? _GEN_9 : _GEN_377; // @[TBE.scala 109:24]
  wire [31:0] _GEN_443 = isAlloc_0 ? _GEN_10 : _GEN_378; // @[TBE.scala 109:24]
  wire [31:0] _GEN_444 = isAlloc_0 ? _GEN_11 : _GEN_379; // @[TBE.scala 109:24]
  wire [31:0] _GEN_445 = isAlloc_0 ? _GEN_12 : _GEN_380; // @[TBE.scala 109:24]
  wire [31:0] _GEN_446 = isAlloc_0 ? _GEN_13 : _GEN_381; // @[TBE.scala 109:24]
  wire [31:0] _GEN_447 = isAlloc_0 ? _GEN_14 : _GEN_382; // @[TBE.scala 109:24]
  wire [31:0] _GEN_448 = isAlloc_0 ? _GEN_15 : _GEN_383; // @[TBE.scala 109:24]
  wire [2:0] _GEN_449 = isAlloc_0 ? _GEN_16 : _GEN_384; // @[TBE.scala 109:24]
  wire [2:0] _GEN_450 = isAlloc_0 ? _GEN_17 : _GEN_385; // @[TBE.scala 109:24]
  wire [2:0] _GEN_451 = isAlloc_0 ? _GEN_18 : _GEN_386; // @[TBE.scala 109:24]
  wire [2:0] _GEN_452 = isAlloc_0 ? _GEN_19 : _GEN_387; // @[TBE.scala 109:24]
  wire [2:0] _GEN_453 = isAlloc_0 ? _GEN_20 : _GEN_388; // @[TBE.scala 109:24]
  wire [2:0] _GEN_454 = isAlloc_0 ? _GEN_21 : _GEN_389; // @[TBE.scala 109:24]
  wire [2:0] _GEN_455 = isAlloc_0 ? _GEN_22 : _GEN_390; // @[TBE.scala 109:24]
  wire [2:0] _GEN_456 = isAlloc_0 ? _GEN_23 : _GEN_391; // @[TBE.scala 109:24]
  wire [2:0] _GEN_457 = isAlloc_0 ? _GEN_24 : _GEN_392; // @[TBE.scala 109:24]
  wire [2:0] _GEN_458 = isAlloc_0 ? _GEN_25 : _GEN_393; // @[TBE.scala 109:24]
  wire [2:0] _GEN_459 = isAlloc_0 ? _GEN_26 : _GEN_394; // @[TBE.scala 109:24]
  wire [2:0] _GEN_460 = isAlloc_0 ? _GEN_27 : _GEN_395; // @[TBE.scala 109:24]
  wire [2:0] _GEN_461 = isAlloc_0 ? _GEN_28 : _GEN_396; // @[TBE.scala 109:24]
  wire [2:0] _GEN_462 = isAlloc_0 ? _GEN_29 : _GEN_397; // @[TBE.scala 109:24]
  wire [2:0] _GEN_463 = isAlloc_0 ? _GEN_30 : _GEN_398; // @[TBE.scala 109:24]
  wire [2:0] _GEN_464 = isAlloc_0 ? _GEN_31 : _GEN_399; // @[TBE.scala 109:24]
  wire [1:0] _GEN_465 = isAlloc_0 ? _GEN_32 : _GEN_400; // @[TBE.scala 109:24]
  wire [1:0] _GEN_466 = isAlloc_0 ? _GEN_33 : _GEN_401; // @[TBE.scala 109:24]
  wire [1:0] _GEN_467 = isAlloc_0 ? _GEN_34 : _GEN_402; // @[TBE.scala 109:24]
  wire [1:0] _GEN_468 = isAlloc_0 ? _GEN_35 : _GEN_403; // @[TBE.scala 109:24]
  wire [1:0] _GEN_469 = isAlloc_0 ? _GEN_36 : _GEN_404; // @[TBE.scala 109:24]
  wire [1:0] _GEN_470 = isAlloc_0 ? _GEN_37 : _GEN_405; // @[TBE.scala 109:24]
  wire [1:0] _GEN_471 = isAlloc_0 ? _GEN_38 : _GEN_406; // @[TBE.scala 109:24]
  wire [1:0] _GEN_472 = isAlloc_0 ? _GEN_39 : _GEN_407; // @[TBE.scala 109:24]
  wire [1:0] _GEN_473 = isAlloc_0 ? _GEN_40 : _GEN_408; // @[TBE.scala 109:24]
  wire [1:0] _GEN_474 = isAlloc_0 ? _GEN_41 : _GEN_409; // @[TBE.scala 109:24]
  wire [1:0] _GEN_475 = isAlloc_0 ? _GEN_42 : _GEN_410; // @[TBE.scala 109:24]
  wire [1:0] _GEN_476 = isAlloc_0 ? _GEN_43 : _GEN_411; // @[TBE.scala 109:24]
  wire [1:0] _GEN_477 = isAlloc_0 ? _GEN_44 : _GEN_412; // @[TBE.scala 109:24]
  wire [1:0] _GEN_478 = isAlloc_0 ? _GEN_45 : _GEN_413; // @[TBE.scala 109:24]
  wire [1:0] _GEN_479 = isAlloc_0 ? _GEN_46 : _GEN_414; // @[TBE.scala 109:24]
  wire [1:0] _GEN_480 = isAlloc_0 ? _GEN_47 : _GEN_415; // @[TBE.scala 109:24]
  wire [31:0] _GEN_481 = isAlloc_0 ? _GEN_48 : _GEN_416; // @[TBE.scala 109:24]
  wire [31:0] _GEN_482 = isAlloc_0 ? _GEN_49 : _GEN_417; // @[TBE.scala 109:24]
  wire [31:0] _GEN_483 = isAlloc_0 ? _GEN_50 : _GEN_418; // @[TBE.scala 109:24]
  wire [31:0] _GEN_484 = isAlloc_0 ? _GEN_51 : _GEN_419; // @[TBE.scala 109:24]
  wire [31:0] _GEN_485 = isAlloc_0 ? _GEN_52 : _GEN_420; // @[TBE.scala 109:24]
  wire [31:0] _GEN_486 = isAlloc_0 ? _GEN_53 : _GEN_421; // @[TBE.scala 109:24]
  wire [31:0] _GEN_487 = isAlloc_0 ? _GEN_54 : _GEN_422; // @[TBE.scala 109:24]
  wire [31:0] _GEN_488 = isAlloc_0 ? _GEN_55 : _GEN_423; // @[TBE.scala 109:24]
  wire [31:0] _GEN_489 = isAlloc_0 ? _GEN_56 : _GEN_424; // @[TBE.scala 109:24]
  wire [31:0] _GEN_490 = isAlloc_0 ? _GEN_57 : _GEN_425; // @[TBE.scala 109:24]
  wire [31:0] _GEN_491 = isAlloc_0 ? _GEN_58 : _GEN_426; // @[TBE.scala 109:24]
  wire [31:0] _GEN_492 = isAlloc_0 ? _GEN_59 : _GEN_427; // @[TBE.scala 109:24]
  wire [31:0] _GEN_493 = isAlloc_0 ? _GEN_60 : _GEN_428; // @[TBE.scala 109:24]
  wire [31:0] _GEN_494 = isAlloc_0 ? _GEN_61 : _GEN_429; // @[TBE.scala 109:24]
  wire [31:0] _GEN_495 = isAlloc_0 ? _GEN_62 : _GEN_430; // @[TBE.scala 109:24]
  wire [31:0] _GEN_496 = isAlloc_0 ? _GEN_63 : _GEN_431; // @[TBE.scala 109:24]
  wire  _GEN_497 = isAlloc_0 ? _GEN_64 : _GEN_352; // @[TBE.scala 109:24]
  wire  _GEN_498 = isAlloc_0 ? _GEN_65 : _GEN_353; // @[TBE.scala 109:24]
  wire  _GEN_499 = isAlloc_0 ? _GEN_66 : _GEN_354; // @[TBE.scala 109:24]
  wire  _GEN_500 = isAlloc_0 ? _GEN_67 : _GEN_355; // @[TBE.scala 109:24]
  wire  _GEN_501 = isAlloc_0 ? _GEN_68 : _GEN_356; // @[TBE.scala 109:24]
  wire  _GEN_502 = isAlloc_0 ? _GEN_69 : _GEN_357; // @[TBE.scala 109:24]
  wire  _GEN_503 = isAlloc_0 ? _GEN_70 : _GEN_358; // @[TBE.scala 109:24]
  wire  _GEN_504 = isAlloc_0 ? _GEN_71 : _GEN_359; // @[TBE.scala 109:24]
  wire  _GEN_505 = isAlloc_0 ? _GEN_72 : _GEN_360; // @[TBE.scala 109:24]
  wire  _GEN_506 = isAlloc_0 ? _GEN_73 : _GEN_361; // @[TBE.scala 109:24]
  wire  _GEN_507 = isAlloc_0 ? _GEN_74 : _GEN_362; // @[TBE.scala 109:24]
  wire  _GEN_508 = isAlloc_0 ? _GEN_75 : _GEN_363; // @[TBE.scala 109:24]
  wire  _GEN_509 = isAlloc_0 ? _GEN_76 : _GEN_364; // @[TBE.scala 109:24]
  wire  _GEN_510 = isAlloc_0 ? _GEN_77 : _GEN_365; // @[TBE.scala 109:24]
  wire  _GEN_511 = isAlloc_0 ? _GEN_78 : _GEN_366; // @[TBE.scala 109:24]
  wire  _GEN_512 = isAlloc_0 ? _GEN_79 : _GEN_367; // @[TBE.scala 109:24]
  wire [31:0] _GEN_514 = 4'h0 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_433; // @[TBE.scala 110:27]
  wire [31:0] _GEN_515 = 4'h1 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_434; // @[TBE.scala 110:27]
  wire [31:0] _GEN_516 = 4'h2 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_435; // @[TBE.scala 110:27]
  wire [31:0] _GEN_517 = 4'h3 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_436; // @[TBE.scala 110:27]
  wire [31:0] _GEN_518 = 4'h4 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_437; // @[TBE.scala 110:27]
  wire [31:0] _GEN_519 = 4'h5 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_438; // @[TBE.scala 110:27]
  wire [31:0] _GEN_520 = 4'h6 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_439; // @[TBE.scala 110:27]
  wire [31:0] _GEN_521 = 4'h7 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_440; // @[TBE.scala 110:27]
  wire [31:0] _GEN_522 = 4'h8 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_441; // @[TBE.scala 110:27]
  wire [31:0] _GEN_523 = 4'h9 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_442; // @[TBE.scala 110:27]
  wire [31:0] _GEN_524 = 4'ha == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_443; // @[TBE.scala 110:27]
  wire [31:0] _GEN_525 = 4'hb == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_444; // @[TBE.scala 110:27]
  wire [31:0] _GEN_526 = 4'hc == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_445; // @[TBE.scala 110:27]
  wire [31:0] _GEN_527 = 4'hd == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_446; // @[TBE.scala 110:27]
  wire [31:0] _GEN_528 = 4'he == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_447; // @[TBE.scala 110:27]
  wire [31:0] _GEN_529 = 4'hf == idxAlloc[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_448; // @[TBE.scala 110:27]
  wire [2:0] _GEN_530 = 4'h0 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_449; // @[TBE.scala 110:27]
  wire [2:0] _GEN_531 = 4'h1 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_450; // @[TBE.scala 110:27]
  wire [2:0] _GEN_532 = 4'h2 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_451; // @[TBE.scala 110:27]
  wire [2:0] _GEN_533 = 4'h3 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_452; // @[TBE.scala 110:27]
  wire [2:0] _GEN_534 = 4'h4 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_453; // @[TBE.scala 110:27]
  wire [2:0] _GEN_535 = 4'h5 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_454; // @[TBE.scala 110:27]
  wire [2:0] _GEN_536 = 4'h6 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_455; // @[TBE.scala 110:27]
  wire [2:0] _GEN_537 = 4'h7 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_456; // @[TBE.scala 110:27]
  wire [2:0] _GEN_538 = 4'h8 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_457; // @[TBE.scala 110:27]
  wire [2:0] _GEN_539 = 4'h9 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_458; // @[TBE.scala 110:27]
  wire [2:0] _GEN_540 = 4'ha == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_459; // @[TBE.scala 110:27]
  wire [2:0] _GEN_541 = 4'hb == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_460; // @[TBE.scala 110:27]
  wire [2:0] _GEN_542 = 4'hc == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_461; // @[TBE.scala 110:27]
  wire [2:0] _GEN_543 = 4'hd == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_462; // @[TBE.scala 110:27]
  wire [2:0] _GEN_544 = 4'he == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_463; // @[TBE.scala 110:27]
  wire [2:0] _GEN_545 = 4'hf == idxAlloc[3:0] ? io_write_1_bits_inputTBE_way : _GEN_464; // @[TBE.scala 110:27]
  wire [1:0] _GEN_546 = 4'h0 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_465; // @[TBE.scala 110:27]
  wire [1:0] _GEN_547 = 4'h1 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_466; // @[TBE.scala 110:27]
  wire [1:0] _GEN_548 = 4'h2 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_467; // @[TBE.scala 110:27]
  wire [1:0] _GEN_549 = 4'h3 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_468; // @[TBE.scala 110:27]
  wire [1:0] _GEN_550 = 4'h4 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_469; // @[TBE.scala 110:27]
  wire [1:0] _GEN_551 = 4'h5 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_470; // @[TBE.scala 110:27]
  wire [1:0] _GEN_552 = 4'h6 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_471; // @[TBE.scala 110:27]
  wire [1:0] _GEN_553 = 4'h7 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_472; // @[TBE.scala 110:27]
  wire [1:0] _GEN_554 = 4'h8 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_473; // @[TBE.scala 110:27]
  wire [1:0] _GEN_555 = 4'h9 == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_474; // @[TBE.scala 110:27]
  wire [1:0] _GEN_556 = 4'ha == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_475; // @[TBE.scala 110:27]
  wire [1:0] _GEN_557 = 4'hb == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_476; // @[TBE.scala 110:27]
  wire [1:0] _GEN_558 = 4'hc == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_477; // @[TBE.scala 110:27]
  wire [1:0] _GEN_559 = 4'hd == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_478; // @[TBE.scala 110:27]
  wire [1:0] _GEN_560 = 4'he == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_479; // @[TBE.scala 110:27]
  wire [1:0] _GEN_561 = 4'hf == idxAlloc[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_480; // @[TBE.scala 110:27]
  wire [31:0] _GEN_562 = 4'h0 == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_481; // @[TBE.scala 111:25]
  wire [31:0] _GEN_563 = 4'h1 == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_482; // @[TBE.scala 111:25]
  wire [31:0] _GEN_564 = 4'h2 == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_483; // @[TBE.scala 111:25]
  wire [31:0] _GEN_565 = 4'h3 == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_484; // @[TBE.scala 111:25]
  wire [31:0] _GEN_566 = 4'h4 == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_485; // @[TBE.scala 111:25]
  wire [31:0] _GEN_567 = 4'h5 == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_486; // @[TBE.scala 111:25]
  wire [31:0] _GEN_568 = 4'h6 == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_487; // @[TBE.scala 111:25]
  wire [31:0] _GEN_569 = 4'h7 == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_488; // @[TBE.scala 111:25]
  wire [31:0] _GEN_570 = 4'h8 == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_489; // @[TBE.scala 111:25]
  wire [31:0] _GEN_571 = 4'h9 == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_490; // @[TBE.scala 111:25]
  wire [31:0] _GEN_572 = 4'ha == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_491; // @[TBE.scala 111:25]
  wire [31:0] _GEN_573 = 4'hb == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_492; // @[TBE.scala 111:25]
  wire [31:0] _GEN_574 = 4'hc == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_493; // @[TBE.scala 111:25]
  wire [31:0] _GEN_575 = 4'hd == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_494; // @[TBE.scala 111:25]
  wire [31:0] _GEN_576 = 4'he == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_495; // @[TBE.scala 111:25]
  wire [31:0] _GEN_577 = 4'hf == idxAlloc[3:0] ? io_write_1_bits_addr[31:0] : _GEN_496; // @[TBE.scala 111:25]
  wire  _GEN_578 = _GEN_4161 | _GEN_497; // @[TBE.scala 112:26]
  wire  _GEN_579 = _GEN_4162 | _GEN_498; // @[TBE.scala 112:26]
  wire  _GEN_580 = _GEN_4163 | _GEN_499; // @[TBE.scala 112:26]
  wire  _GEN_581 = _GEN_4164 | _GEN_500; // @[TBE.scala 112:26]
  wire  _GEN_582 = _GEN_4165 | _GEN_501; // @[TBE.scala 112:26]
  wire  _GEN_583 = _GEN_4166 | _GEN_502; // @[TBE.scala 112:26]
  wire  _GEN_584 = _GEN_4167 | _GEN_503; // @[TBE.scala 112:26]
  wire  _GEN_585 = _GEN_4168 | _GEN_504; // @[TBE.scala 112:26]
  wire  _GEN_586 = _GEN_4169 | _GEN_505; // @[TBE.scala 112:26]
  wire  _GEN_587 = _GEN_4170 | _GEN_506; // @[TBE.scala 112:26]
  wire  _GEN_588 = _GEN_4171 | _GEN_507; // @[TBE.scala 112:26]
  wire  _GEN_589 = _GEN_4172 | _GEN_508; // @[TBE.scala 112:26]
  wire  _GEN_590 = _GEN_4173 | _GEN_509; // @[TBE.scala 112:26]
  wire  _GEN_591 = _GEN_4174 | _GEN_510; // @[TBE.scala 112:26]
  wire  _GEN_592 = _GEN_4175 | _GEN_511; // @[TBE.scala 112:26]
  wire  _GEN_593 = _GEN_4176 | _GEN_512; // @[TBE.scala 112:26]
  wire  _T_271 = io_write_1_bits_command == 2'h2; // @[TBE.scala 137:46]
  wire  isDealloc_1 = _T_271 & io_write_1_valid; // @[TBE.scala 137:58]
  wire  _T_111 = isDealloc_1 & finder_1_io_value_valid; // @[TBE.scala 114:31]
  wire [4:0] idxUpdate_1 = {{1'd0}, finder_1_io_value_bits}; // @[TBE.scala 73:23 TBE.scala 104:18]
  wire  _GEN_594 = 4'h0 == idxUpdate_1[3:0] ? 1'h0 : _GEN_497; // @[TBE.scala 115:30]
  wire  _GEN_595 = 4'h1 == idxUpdate_1[3:0] ? 1'h0 : _GEN_498; // @[TBE.scala 115:30]
  wire  _GEN_596 = 4'h2 == idxUpdate_1[3:0] ? 1'h0 : _GEN_499; // @[TBE.scala 115:30]
  wire  _GEN_597 = 4'h3 == idxUpdate_1[3:0] ? 1'h0 : _GEN_500; // @[TBE.scala 115:30]
  wire  _GEN_598 = 4'h4 == idxUpdate_1[3:0] ? 1'h0 : _GEN_501; // @[TBE.scala 115:30]
  wire  _GEN_599 = 4'h5 == idxUpdate_1[3:0] ? 1'h0 : _GEN_502; // @[TBE.scala 115:30]
  wire  _GEN_600 = 4'h6 == idxUpdate_1[3:0] ? 1'h0 : _GEN_503; // @[TBE.scala 115:30]
  wire  _GEN_601 = 4'h7 == idxUpdate_1[3:0] ? 1'h0 : _GEN_504; // @[TBE.scala 115:30]
  wire  _GEN_602 = 4'h8 == idxUpdate_1[3:0] ? 1'h0 : _GEN_505; // @[TBE.scala 115:30]
  wire  _GEN_603 = 4'h9 == idxUpdate_1[3:0] ? 1'h0 : _GEN_506; // @[TBE.scala 115:30]
  wire  _GEN_604 = 4'ha == idxUpdate_1[3:0] ? 1'h0 : _GEN_507; // @[TBE.scala 115:30]
  wire  _GEN_605 = 4'hb == idxUpdate_1[3:0] ? 1'h0 : _GEN_508; // @[TBE.scala 115:30]
  wire  _GEN_606 = 4'hc == idxUpdate_1[3:0] ? 1'h0 : _GEN_509; // @[TBE.scala 115:30]
  wire  _GEN_607 = 4'hd == idxUpdate_1[3:0] ? 1'h0 : _GEN_510; // @[TBE.scala 115:30]
  wire  _GEN_608 = 4'he == idxUpdate_1[3:0] ? 1'h0 : _GEN_511; // @[TBE.scala 115:30]
  wire  _GEN_609 = 4'hf == idxUpdate_1[3:0] ? 1'h0 : _GEN_512; // @[TBE.scala 115:30]
  wire [31:0] _GEN_610 = 4'h0 == idxUpdate_1[3:0] ? 32'h0 : _GEN_433; // @[TBE.scala 116:31]
  wire [31:0] _GEN_611 = 4'h1 == idxUpdate_1[3:0] ? 32'h0 : _GEN_434; // @[TBE.scala 116:31]
  wire [31:0] _GEN_612 = 4'h2 == idxUpdate_1[3:0] ? 32'h0 : _GEN_435; // @[TBE.scala 116:31]
  wire [31:0] _GEN_613 = 4'h3 == idxUpdate_1[3:0] ? 32'h0 : _GEN_436; // @[TBE.scala 116:31]
  wire [31:0] _GEN_614 = 4'h4 == idxUpdate_1[3:0] ? 32'h0 : _GEN_437; // @[TBE.scala 116:31]
  wire [31:0] _GEN_615 = 4'h5 == idxUpdate_1[3:0] ? 32'h0 : _GEN_438; // @[TBE.scala 116:31]
  wire [31:0] _GEN_616 = 4'h6 == idxUpdate_1[3:0] ? 32'h0 : _GEN_439; // @[TBE.scala 116:31]
  wire [31:0] _GEN_617 = 4'h7 == idxUpdate_1[3:0] ? 32'h0 : _GEN_440; // @[TBE.scala 116:31]
  wire [31:0] _GEN_618 = 4'h8 == idxUpdate_1[3:0] ? 32'h0 : _GEN_441; // @[TBE.scala 116:31]
  wire [31:0] _GEN_619 = 4'h9 == idxUpdate_1[3:0] ? 32'h0 : _GEN_442; // @[TBE.scala 116:31]
  wire [31:0] _GEN_620 = 4'ha == idxUpdate_1[3:0] ? 32'h0 : _GEN_443; // @[TBE.scala 116:31]
  wire [31:0] _GEN_621 = 4'hb == idxUpdate_1[3:0] ? 32'h0 : _GEN_444; // @[TBE.scala 116:31]
  wire [31:0] _GEN_622 = 4'hc == idxUpdate_1[3:0] ? 32'h0 : _GEN_445; // @[TBE.scala 116:31]
  wire [31:0] _GEN_623 = 4'hd == idxUpdate_1[3:0] ? 32'h0 : _GEN_446; // @[TBE.scala 116:31]
  wire [31:0] _GEN_624 = 4'he == idxUpdate_1[3:0] ? 32'h0 : _GEN_447; // @[TBE.scala 116:31]
  wire [31:0] _GEN_625 = 4'hf == idxUpdate_1[3:0] ? 32'h0 : _GEN_448; // @[TBE.scala 116:31]
  wire [2:0] _GEN_626 = 4'h0 == idxUpdate_1[3:0] ? 3'h2 : _GEN_449; // @[TBE.scala 116:31]
  wire [2:0] _GEN_627 = 4'h1 == idxUpdate_1[3:0] ? 3'h2 : _GEN_450; // @[TBE.scala 116:31]
  wire [2:0] _GEN_628 = 4'h2 == idxUpdate_1[3:0] ? 3'h2 : _GEN_451; // @[TBE.scala 116:31]
  wire [2:0] _GEN_629 = 4'h3 == idxUpdate_1[3:0] ? 3'h2 : _GEN_452; // @[TBE.scala 116:31]
  wire [2:0] _GEN_630 = 4'h4 == idxUpdate_1[3:0] ? 3'h2 : _GEN_453; // @[TBE.scala 116:31]
  wire [2:0] _GEN_631 = 4'h5 == idxUpdate_1[3:0] ? 3'h2 : _GEN_454; // @[TBE.scala 116:31]
  wire [2:0] _GEN_632 = 4'h6 == idxUpdate_1[3:0] ? 3'h2 : _GEN_455; // @[TBE.scala 116:31]
  wire [2:0] _GEN_633 = 4'h7 == idxUpdate_1[3:0] ? 3'h2 : _GEN_456; // @[TBE.scala 116:31]
  wire [2:0] _GEN_634 = 4'h8 == idxUpdate_1[3:0] ? 3'h2 : _GEN_457; // @[TBE.scala 116:31]
  wire [2:0] _GEN_635 = 4'h9 == idxUpdate_1[3:0] ? 3'h2 : _GEN_458; // @[TBE.scala 116:31]
  wire [2:0] _GEN_636 = 4'ha == idxUpdate_1[3:0] ? 3'h2 : _GEN_459; // @[TBE.scala 116:31]
  wire [2:0] _GEN_637 = 4'hb == idxUpdate_1[3:0] ? 3'h2 : _GEN_460; // @[TBE.scala 116:31]
  wire [2:0] _GEN_638 = 4'hc == idxUpdate_1[3:0] ? 3'h2 : _GEN_461; // @[TBE.scala 116:31]
  wire [2:0] _GEN_639 = 4'hd == idxUpdate_1[3:0] ? 3'h2 : _GEN_462; // @[TBE.scala 116:31]
  wire [2:0] _GEN_640 = 4'he == idxUpdate_1[3:0] ? 3'h2 : _GEN_463; // @[TBE.scala 116:31]
  wire [2:0] _GEN_641 = 4'hf == idxUpdate_1[3:0] ? 3'h2 : _GEN_464; // @[TBE.scala 116:31]
  wire [1:0] _GEN_642 = 4'h0 == idxUpdate_1[3:0] ? 2'h0 : _GEN_465; // @[TBE.scala 116:31]
  wire [1:0] _GEN_643 = 4'h1 == idxUpdate_1[3:0] ? 2'h0 : _GEN_466; // @[TBE.scala 116:31]
  wire [1:0] _GEN_644 = 4'h2 == idxUpdate_1[3:0] ? 2'h0 : _GEN_467; // @[TBE.scala 116:31]
  wire [1:0] _GEN_645 = 4'h3 == idxUpdate_1[3:0] ? 2'h0 : _GEN_468; // @[TBE.scala 116:31]
  wire [1:0] _GEN_646 = 4'h4 == idxUpdate_1[3:0] ? 2'h0 : _GEN_469; // @[TBE.scala 116:31]
  wire [1:0] _GEN_647 = 4'h5 == idxUpdate_1[3:0] ? 2'h0 : _GEN_470; // @[TBE.scala 116:31]
  wire [1:0] _GEN_648 = 4'h6 == idxUpdate_1[3:0] ? 2'h0 : _GEN_471; // @[TBE.scala 116:31]
  wire [1:0] _GEN_649 = 4'h7 == idxUpdate_1[3:0] ? 2'h0 : _GEN_472; // @[TBE.scala 116:31]
  wire [1:0] _GEN_650 = 4'h8 == idxUpdate_1[3:0] ? 2'h0 : _GEN_473; // @[TBE.scala 116:31]
  wire [1:0] _GEN_651 = 4'h9 == idxUpdate_1[3:0] ? 2'h0 : _GEN_474; // @[TBE.scala 116:31]
  wire [1:0] _GEN_652 = 4'ha == idxUpdate_1[3:0] ? 2'h0 : _GEN_475; // @[TBE.scala 116:31]
  wire [1:0] _GEN_653 = 4'hb == idxUpdate_1[3:0] ? 2'h0 : _GEN_476; // @[TBE.scala 116:31]
  wire [1:0] _GEN_654 = 4'hc == idxUpdate_1[3:0] ? 2'h0 : _GEN_477; // @[TBE.scala 116:31]
  wire [1:0] _GEN_655 = 4'hd == idxUpdate_1[3:0] ? 2'h0 : _GEN_478; // @[TBE.scala 116:31]
  wire [1:0] _GEN_656 = 4'he == idxUpdate_1[3:0] ? 2'h0 : _GEN_479; // @[TBE.scala 116:31]
  wire [1:0] _GEN_657 = 4'hf == idxUpdate_1[3:0] ? 2'h0 : _GEN_480; // @[TBE.scala 116:31]
  wire [31:0] _GEN_658 = 4'h0 == idxUpdate_1[3:0] ? 32'h0 : _GEN_481; // @[TBE.scala 117:29]
  wire [31:0] _GEN_659 = 4'h1 == idxUpdate_1[3:0] ? 32'h0 : _GEN_482; // @[TBE.scala 117:29]
  wire [31:0] _GEN_660 = 4'h2 == idxUpdate_1[3:0] ? 32'h0 : _GEN_483; // @[TBE.scala 117:29]
  wire [31:0] _GEN_661 = 4'h3 == idxUpdate_1[3:0] ? 32'h0 : _GEN_484; // @[TBE.scala 117:29]
  wire [31:0] _GEN_662 = 4'h4 == idxUpdate_1[3:0] ? 32'h0 : _GEN_485; // @[TBE.scala 117:29]
  wire [31:0] _GEN_663 = 4'h5 == idxUpdate_1[3:0] ? 32'h0 : _GEN_486; // @[TBE.scala 117:29]
  wire [31:0] _GEN_664 = 4'h6 == idxUpdate_1[3:0] ? 32'h0 : _GEN_487; // @[TBE.scala 117:29]
  wire [31:0] _GEN_665 = 4'h7 == idxUpdate_1[3:0] ? 32'h0 : _GEN_488; // @[TBE.scala 117:29]
  wire [31:0] _GEN_666 = 4'h8 == idxUpdate_1[3:0] ? 32'h0 : _GEN_489; // @[TBE.scala 117:29]
  wire [31:0] _GEN_667 = 4'h9 == idxUpdate_1[3:0] ? 32'h0 : _GEN_490; // @[TBE.scala 117:29]
  wire [31:0] _GEN_668 = 4'ha == idxUpdate_1[3:0] ? 32'h0 : _GEN_491; // @[TBE.scala 117:29]
  wire [31:0] _GEN_669 = 4'hb == idxUpdate_1[3:0] ? 32'h0 : _GEN_492; // @[TBE.scala 117:29]
  wire [31:0] _GEN_670 = 4'hc == idxUpdate_1[3:0] ? 32'h0 : _GEN_493; // @[TBE.scala 117:29]
  wire [31:0] _GEN_671 = 4'hd == idxUpdate_1[3:0] ? 32'h0 : _GEN_494; // @[TBE.scala 117:29]
  wire [31:0] _GEN_672 = 4'he == idxUpdate_1[3:0] ? 32'h0 : _GEN_495; // @[TBE.scala 117:29]
  wire [31:0] _GEN_673 = 4'hf == idxUpdate_1[3:0] ? 32'h0 : _GEN_496; // @[TBE.scala 117:29]
  wire  _T_273 = io_write_1_bits_command == 2'h3; // @[TBE.scala 138:44]
  wire  isWrite_1 = _T_273 & io_write_1_valid; // @[TBE.scala 138:55]
  wire  _T_119 = isWrite_1 & finder_1_io_value_valid; // @[TBE.scala 119:29]
  wire  _T_120 = ~io_write_1_bits_mask; // @[TBE.scala 120:35]
  wire [31:0] _GEN_674 = 4'h0 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_433; // @[TBE.scala 121:63]
  wire [31:0] _GEN_675 = 4'h1 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_434; // @[TBE.scala 121:63]
  wire [31:0] _GEN_676 = 4'h2 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_435; // @[TBE.scala 121:63]
  wire [31:0] _GEN_677 = 4'h3 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_436; // @[TBE.scala 121:63]
  wire [31:0] _GEN_678 = 4'h4 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_437; // @[TBE.scala 121:63]
  wire [31:0] _GEN_679 = 4'h5 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_438; // @[TBE.scala 121:63]
  wire [31:0] _GEN_680 = 4'h6 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_439; // @[TBE.scala 121:63]
  wire [31:0] _GEN_681 = 4'h7 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_440; // @[TBE.scala 121:63]
  wire [31:0] _GEN_682 = 4'h8 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_441; // @[TBE.scala 121:63]
  wire [31:0] _GEN_683 = 4'h9 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_442; // @[TBE.scala 121:63]
  wire [31:0] _GEN_684 = 4'ha == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_443; // @[TBE.scala 121:63]
  wire [31:0] _GEN_685 = 4'hb == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_444; // @[TBE.scala 121:63]
  wire [31:0] _GEN_686 = 4'hc == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_445; // @[TBE.scala 121:63]
  wire [31:0] _GEN_687 = 4'hd == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_446; // @[TBE.scala 121:63]
  wire [31:0] _GEN_688 = 4'he == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_447; // @[TBE.scala 121:63]
  wire [31:0] _GEN_689 = 4'hf == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_fields_0 : _GEN_448; // @[TBE.scala 121:63]
  wire [31:0] _GEN_695 = 4'h1 == idxUpdate_1[3:0] ? TBEMemory_1_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 122:15]
  wire [31:0] _GEN_698 = 4'h2 == idxUpdate_1[3:0] ? TBEMemory_2_fields_0 : _GEN_695; // @[TBE.scala 122:15]
  wire [31:0] _GEN_701 = 4'h3 == idxUpdate_1[3:0] ? TBEMemory_3_fields_0 : _GEN_698; // @[TBE.scala 122:15]
  wire [31:0] _GEN_704 = 4'h4 == idxUpdate_1[3:0] ? TBEMemory_4_fields_0 : _GEN_701; // @[TBE.scala 122:15]
  wire [31:0] _GEN_707 = 4'h5 == idxUpdate_1[3:0] ? TBEMemory_5_fields_0 : _GEN_704; // @[TBE.scala 122:15]
  wire [31:0] _GEN_710 = 4'h6 == idxUpdate_1[3:0] ? TBEMemory_6_fields_0 : _GEN_707; // @[TBE.scala 122:15]
  wire [31:0] _GEN_713 = 4'h7 == idxUpdate_1[3:0] ? TBEMemory_7_fields_0 : _GEN_710; // @[TBE.scala 122:15]
  wire [31:0] _GEN_716 = 4'h8 == idxUpdate_1[3:0] ? TBEMemory_8_fields_0 : _GEN_713; // @[TBE.scala 122:15]
  wire [31:0] _GEN_719 = 4'h9 == idxUpdate_1[3:0] ? TBEMemory_9_fields_0 : _GEN_716; // @[TBE.scala 122:15]
  wire [31:0] _GEN_722 = 4'ha == idxUpdate_1[3:0] ? TBEMemory_10_fields_0 : _GEN_719; // @[TBE.scala 122:15]
  wire [31:0] _GEN_725 = 4'hb == idxUpdate_1[3:0] ? TBEMemory_11_fields_0 : _GEN_722; // @[TBE.scala 122:15]
  wire [31:0] _GEN_728 = 4'hc == idxUpdate_1[3:0] ? TBEMemory_12_fields_0 : _GEN_725; // @[TBE.scala 122:15]
  wire [31:0] _GEN_731 = 4'hd == idxUpdate_1[3:0] ? TBEMemory_13_fields_0 : _GEN_728; // @[TBE.scala 122:15]
  wire [31:0] _GEN_734 = 4'he == idxUpdate_1[3:0] ? TBEMemory_14_fields_0 : _GEN_731; // @[TBE.scala 122:15]
  wire [31:0] _GEN_737 = 4'hf == idxUpdate_1[3:0] ? TBEMemory_15_fields_0 : _GEN_734; // @[TBE.scala 122:15]
  wire [2:0] _GEN_738 = 4'h0 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_449; // @[TBE.scala 124:37]
  wire [2:0] _GEN_739 = 4'h1 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_450; // @[TBE.scala 124:37]
  wire [2:0] _GEN_740 = 4'h2 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_451; // @[TBE.scala 124:37]
  wire [2:0] _GEN_741 = 4'h3 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_452; // @[TBE.scala 124:37]
  wire [2:0] _GEN_742 = 4'h4 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_453; // @[TBE.scala 124:37]
  wire [2:0] _GEN_743 = 4'h5 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_454; // @[TBE.scala 124:37]
  wire [2:0] _GEN_744 = 4'h6 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_455; // @[TBE.scala 124:37]
  wire [2:0] _GEN_745 = 4'h7 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_456; // @[TBE.scala 124:37]
  wire [2:0] _GEN_746 = 4'h8 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_457; // @[TBE.scala 124:37]
  wire [2:0] _GEN_747 = 4'h9 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_458; // @[TBE.scala 124:37]
  wire [2:0] _GEN_748 = 4'ha == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_459; // @[TBE.scala 124:37]
  wire [2:0] _GEN_749 = 4'hb == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_460; // @[TBE.scala 124:37]
  wire [2:0] _GEN_750 = 4'hc == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_461; // @[TBE.scala 124:37]
  wire [2:0] _GEN_751 = 4'hd == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_462; // @[TBE.scala 124:37]
  wire [2:0] _GEN_752 = 4'he == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_463; // @[TBE.scala 124:37]
  wire [2:0] _GEN_753 = 4'hf == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_way : _GEN_464; // @[TBE.scala 124:37]
  wire [1:0] _GEN_754 = 4'h0 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_465; // @[TBE.scala 125:39]
  wire [1:0] _GEN_755 = 4'h1 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_466; // @[TBE.scala 125:39]
  wire [1:0] _GEN_756 = 4'h2 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_467; // @[TBE.scala 125:39]
  wire [1:0] _GEN_757 = 4'h3 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_468; // @[TBE.scala 125:39]
  wire [1:0] _GEN_758 = 4'h4 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_469; // @[TBE.scala 125:39]
  wire [1:0] _GEN_759 = 4'h5 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_470; // @[TBE.scala 125:39]
  wire [1:0] _GEN_760 = 4'h6 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_471; // @[TBE.scala 125:39]
  wire [1:0] _GEN_761 = 4'h7 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_472; // @[TBE.scala 125:39]
  wire [1:0] _GEN_762 = 4'h8 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_473; // @[TBE.scala 125:39]
  wire [1:0] _GEN_763 = 4'h9 == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_474; // @[TBE.scala 125:39]
  wire [1:0] _GEN_764 = 4'ha == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_475; // @[TBE.scala 125:39]
  wire [1:0] _GEN_765 = 4'hb == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_476; // @[TBE.scala 125:39]
  wire [1:0] _GEN_766 = 4'hc == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_477; // @[TBE.scala 125:39]
  wire [1:0] _GEN_767 = 4'hd == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_478; // @[TBE.scala 125:39]
  wire [1:0] _GEN_768 = 4'he == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_479; // @[TBE.scala 125:39]
  wire [1:0] _GEN_769 = 4'hf == idxUpdate_1[3:0] ? io_write_1_bits_inputTBE_state_state : _GEN_480; // @[TBE.scala 125:39]
  wire [31:0] _GEN_770 = _T_120 ? _GEN_674 : _GEN_433; // @[TBE.scala 120:53]
  wire [31:0] _GEN_771 = _T_120 ? _GEN_675 : _GEN_434; // @[TBE.scala 120:53]
  wire [31:0] _GEN_772 = _T_120 ? _GEN_676 : _GEN_435; // @[TBE.scala 120:53]
  wire [31:0] _GEN_773 = _T_120 ? _GEN_677 : _GEN_436; // @[TBE.scala 120:53]
  wire [31:0] _GEN_774 = _T_120 ? _GEN_678 : _GEN_437; // @[TBE.scala 120:53]
  wire [31:0] _GEN_775 = _T_120 ? _GEN_679 : _GEN_438; // @[TBE.scala 120:53]
  wire [31:0] _GEN_776 = _T_120 ? _GEN_680 : _GEN_439; // @[TBE.scala 120:53]
  wire [31:0] _GEN_777 = _T_120 ? _GEN_681 : _GEN_440; // @[TBE.scala 120:53]
  wire [31:0] _GEN_778 = _T_120 ? _GEN_682 : _GEN_441; // @[TBE.scala 120:53]
  wire [31:0] _GEN_779 = _T_120 ? _GEN_683 : _GEN_442; // @[TBE.scala 120:53]
  wire [31:0] _GEN_780 = _T_120 ? _GEN_684 : _GEN_443; // @[TBE.scala 120:53]
  wire [31:0] _GEN_781 = _T_120 ? _GEN_685 : _GEN_444; // @[TBE.scala 120:53]
  wire [31:0] _GEN_782 = _T_120 ? _GEN_686 : _GEN_445; // @[TBE.scala 120:53]
  wire [31:0] _GEN_783 = _T_120 ? _GEN_687 : _GEN_446; // @[TBE.scala 120:53]
  wire [31:0] _GEN_784 = _T_120 ? _GEN_688 : _GEN_447; // @[TBE.scala 120:53]
  wire [31:0] _GEN_785 = _T_120 ? _GEN_689 : _GEN_448; // @[TBE.scala 120:53]
  wire [2:0] _GEN_786 = _T_120 ? _GEN_449 : _GEN_738; // @[TBE.scala 120:53]
  wire [2:0] _GEN_787 = _T_120 ? _GEN_450 : _GEN_739; // @[TBE.scala 120:53]
  wire [2:0] _GEN_788 = _T_120 ? _GEN_451 : _GEN_740; // @[TBE.scala 120:53]
  wire [2:0] _GEN_789 = _T_120 ? _GEN_452 : _GEN_741; // @[TBE.scala 120:53]
  wire [2:0] _GEN_790 = _T_120 ? _GEN_453 : _GEN_742; // @[TBE.scala 120:53]
  wire [2:0] _GEN_791 = _T_120 ? _GEN_454 : _GEN_743; // @[TBE.scala 120:53]
  wire [2:0] _GEN_792 = _T_120 ? _GEN_455 : _GEN_744; // @[TBE.scala 120:53]
  wire [2:0] _GEN_793 = _T_120 ? _GEN_456 : _GEN_745; // @[TBE.scala 120:53]
  wire [2:0] _GEN_794 = _T_120 ? _GEN_457 : _GEN_746; // @[TBE.scala 120:53]
  wire [2:0] _GEN_795 = _T_120 ? _GEN_458 : _GEN_747; // @[TBE.scala 120:53]
  wire [2:0] _GEN_796 = _T_120 ? _GEN_459 : _GEN_748; // @[TBE.scala 120:53]
  wire [2:0] _GEN_797 = _T_120 ? _GEN_460 : _GEN_749; // @[TBE.scala 120:53]
  wire [2:0] _GEN_798 = _T_120 ? _GEN_461 : _GEN_750; // @[TBE.scala 120:53]
  wire [2:0] _GEN_799 = _T_120 ? _GEN_462 : _GEN_751; // @[TBE.scala 120:53]
  wire [2:0] _GEN_800 = _T_120 ? _GEN_463 : _GEN_752; // @[TBE.scala 120:53]
  wire [2:0] _GEN_801 = _T_120 ? _GEN_464 : _GEN_753; // @[TBE.scala 120:53]
  wire [1:0] _GEN_802 = _T_120 ? _GEN_465 : _GEN_754; // @[TBE.scala 120:53]
  wire [1:0] _GEN_803 = _T_120 ? _GEN_466 : _GEN_755; // @[TBE.scala 120:53]
  wire [1:0] _GEN_804 = _T_120 ? _GEN_467 : _GEN_756; // @[TBE.scala 120:53]
  wire [1:0] _GEN_805 = _T_120 ? _GEN_468 : _GEN_757; // @[TBE.scala 120:53]
  wire [1:0] _GEN_806 = _T_120 ? _GEN_469 : _GEN_758; // @[TBE.scala 120:53]
  wire [1:0] _GEN_807 = _T_120 ? _GEN_470 : _GEN_759; // @[TBE.scala 120:53]
  wire [1:0] _GEN_808 = _T_120 ? _GEN_471 : _GEN_760; // @[TBE.scala 120:53]
  wire [1:0] _GEN_809 = _T_120 ? _GEN_472 : _GEN_761; // @[TBE.scala 120:53]
  wire [1:0] _GEN_810 = _T_120 ? _GEN_473 : _GEN_762; // @[TBE.scala 120:53]
  wire [1:0] _GEN_811 = _T_120 ? _GEN_474 : _GEN_763; // @[TBE.scala 120:53]
  wire [1:0] _GEN_812 = _T_120 ? _GEN_475 : _GEN_764; // @[TBE.scala 120:53]
  wire [1:0] _GEN_813 = _T_120 ? _GEN_476 : _GEN_765; // @[TBE.scala 120:53]
  wire [1:0] _GEN_814 = _T_120 ? _GEN_477 : _GEN_766; // @[TBE.scala 120:53]
  wire [1:0] _GEN_815 = _T_120 ? _GEN_478 : _GEN_767; // @[TBE.scala 120:53]
  wire [1:0] _GEN_816 = _T_120 ? _GEN_479 : _GEN_768; // @[TBE.scala 120:53]
  wire [1:0] _GEN_817 = _T_120 ? _GEN_480 : _GEN_769; // @[TBE.scala 120:53]
  wire [31:0] _GEN_818 = _T_119 ? _GEN_770 : _GEN_433; // @[TBE.scala 119:57]
  wire [31:0] _GEN_819 = _T_119 ? _GEN_771 : _GEN_434; // @[TBE.scala 119:57]
  wire [31:0] _GEN_820 = _T_119 ? _GEN_772 : _GEN_435; // @[TBE.scala 119:57]
  wire [31:0] _GEN_821 = _T_119 ? _GEN_773 : _GEN_436; // @[TBE.scala 119:57]
  wire [31:0] _GEN_822 = _T_119 ? _GEN_774 : _GEN_437; // @[TBE.scala 119:57]
  wire [31:0] _GEN_823 = _T_119 ? _GEN_775 : _GEN_438; // @[TBE.scala 119:57]
  wire [31:0] _GEN_824 = _T_119 ? _GEN_776 : _GEN_439; // @[TBE.scala 119:57]
  wire [31:0] _GEN_825 = _T_119 ? _GEN_777 : _GEN_440; // @[TBE.scala 119:57]
  wire [31:0] _GEN_826 = _T_119 ? _GEN_778 : _GEN_441; // @[TBE.scala 119:57]
  wire [31:0] _GEN_827 = _T_119 ? _GEN_779 : _GEN_442; // @[TBE.scala 119:57]
  wire [31:0] _GEN_828 = _T_119 ? _GEN_780 : _GEN_443; // @[TBE.scala 119:57]
  wire [31:0] _GEN_829 = _T_119 ? _GEN_781 : _GEN_444; // @[TBE.scala 119:57]
  wire [31:0] _GEN_830 = _T_119 ? _GEN_782 : _GEN_445; // @[TBE.scala 119:57]
  wire [31:0] _GEN_831 = _T_119 ? _GEN_783 : _GEN_446; // @[TBE.scala 119:57]
  wire [31:0] _GEN_832 = _T_119 ? _GEN_784 : _GEN_447; // @[TBE.scala 119:57]
  wire [31:0] _GEN_833 = _T_119 ? _GEN_785 : _GEN_448; // @[TBE.scala 119:57]
  wire [2:0] _GEN_834 = _T_119 ? _GEN_786 : _GEN_449; // @[TBE.scala 119:57]
  wire [2:0] _GEN_835 = _T_119 ? _GEN_787 : _GEN_450; // @[TBE.scala 119:57]
  wire [2:0] _GEN_836 = _T_119 ? _GEN_788 : _GEN_451; // @[TBE.scala 119:57]
  wire [2:0] _GEN_837 = _T_119 ? _GEN_789 : _GEN_452; // @[TBE.scala 119:57]
  wire [2:0] _GEN_838 = _T_119 ? _GEN_790 : _GEN_453; // @[TBE.scala 119:57]
  wire [2:0] _GEN_839 = _T_119 ? _GEN_791 : _GEN_454; // @[TBE.scala 119:57]
  wire [2:0] _GEN_840 = _T_119 ? _GEN_792 : _GEN_455; // @[TBE.scala 119:57]
  wire [2:0] _GEN_841 = _T_119 ? _GEN_793 : _GEN_456; // @[TBE.scala 119:57]
  wire [2:0] _GEN_842 = _T_119 ? _GEN_794 : _GEN_457; // @[TBE.scala 119:57]
  wire [2:0] _GEN_843 = _T_119 ? _GEN_795 : _GEN_458; // @[TBE.scala 119:57]
  wire [2:0] _GEN_844 = _T_119 ? _GEN_796 : _GEN_459; // @[TBE.scala 119:57]
  wire [2:0] _GEN_845 = _T_119 ? _GEN_797 : _GEN_460; // @[TBE.scala 119:57]
  wire [2:0] _GEN_846 = _T_119 ? _GEN_798 : _GEN_461; // @[TBE.scala 119:57]
  wire [2:0] _GEN_847 = _T_119 ? _GEN_799 : _GEN_462; // @[TBE.scala 119:57]
  wire [2:0] _GEN_848 = _T_119 ? _GEN_800 : _GEN_463; // @[TBE.scala 119:57]
  wire [2:0] _GEN_849 = _T_119 ? _GEN_801 : _GEN_464; // @[TBE.scala 119:57]
  wire [1:0] _GEN_850 = _T_119 ? _GEN_802 : _GEN_465; // @[TBE.scala 119:57]
  wire [1:0] _GEN_851 = _T_119 ? _GEN_803 : _GEN_466; // @[TBE.scala 119:57]
  wire [1:0] _GEN_852 = _T_119 ? _GEN_804 : _GEN_467; // @[TBE.scala 119:57]
  wire [1:0] _GEN_853 = _T_119 ? _GEN_805 : _GEN_468; // @[TBE.scala 119:57]
  wire [1:0] _GEN_854 = _T_119 ? _GEN_806 : _GEN_469; // @[TBE.scala 119:57]
  wire [1:0] _GEN_855 = _T_119 ? _GEN_807 : _GEN_470; // @[TBE.scala 119:57]
  wire [1:0] _GEN_856 = _T_119 ? _GEN_808 : _GEN_471; // @[TBE.scala 119:57]
  wire [1:0] _GEN_857 = _T_119 ? _GEN_809 : _GEN_472; // @[TBE.scala 119:57]
  wire [1:0] _GEN_858 = _T_119 ? _GEN_810 : _GEN_473; // @[TBE.scala 119:57]
  wire [1:0] _GEN_859 = _T_119 ? _GEN_811 : _GEN_474; // @[TBE.scala 119:57]
  wire [1:0] _GEN_860 = _T_119 ? _GEN_812 : _GEN_475; // @[TBE.scala 119:57]
  wire [1:0] _GEN_861 = _T_119 ? _GEN_813 : _GEN_476; // @[TBE.scala 119:57]
  wire [1:0] _GEN_862 = _T_119 ? _GEN_814 : _GEN_477; // @[TBE.scala 119:57]
  wire [1:0] _GEN_863 = _T_119 ? _GEN_815 : _GEN_478; // @[TBE.scala 119:57]
  wire [1:0] _GEN_864 = _T_119 ? _GEN_816 : _GEN_479; // @[TBE.scala 119:57]
  wire [1:0] _GEN_865 = _T_119 ? _GEN_817 : _GEN_480; // @[TBE.scala 119:57]
  wire  _GEN_866 = _T_111 ? _GEN_594 : _GEN_497; // @[TBE.scala 114:59]
  wire  _GEN_867 = _T_111 ? _GEN_595 : _GEN_498; // @[TBE.scala 114:59]
  wire  _GEN_868 = _T_111 ? _GEN_596 : _GEN_499; // @[TBE.scala 114:59]
  wire  _GEN_869 = _T_111 ? _GEN_597 : _GEN_500; // @[TBE.scala 114:59]
  wire  _GEN_870 = _T_111 ? _GEN_598 : _GEN_501; // @[TBE.scala 114:59]
  wire  _GEN_871 = _T_111 ? _GEN_599 : _GEN_502; // @[TBE.scala 114:59]
  wire  _GEN_872 = _T_111 ? _GEN_600 : _GEN_503; // @[TBE.scala 114:59]
  wire  _GEN_873 = _T_111 ? _GEN_601 : _GEN_504; // @[TBE.scala 114:59]
  wire  _GEN_874 = _T_111 ? _GEN_602 : _GEN_505; // @[TBE.scala 114:59]
  wire  _GEN_875 = _T_111 ? _GEN_603 : _GEN_506; // @[TBE.scala 114:59]
  wire  _GEN_876 = _T_111 ? _GEN_604 : _GEN_507; // @[TBE.scala 114:59]
  wire  _GEN_877 = _T_111 ? _GEN_605 : _GEN_508; // @[TBE.scala 114:59]
  wire  _GEN_878 = _T_111 ? _GEN_606 : _GEN_509; // @[TBE.scala 114:59]
  wire  _GEN_879 = _T_111 ? _GEN_607 : _GEN_510; // @[TBE.scala 114:59]
  wire  _GEN_880 = _T_111 ? _GEN_608 : _GEN_511; // @[TBE.scala 114:59]
  wire  _GEN_881 = _T_111 ? _GEN_609 : _GEN_512; // @[TBE.scala 114:59]
  wire [31:0] _GEN_882 = _T_111 ? _GEN_610 : _GEN_818; // @[TBE.scala 114:59]
  wire [31:0] _GEN_883 = _T_111 ? _GEN_611 : _GEN_819; // @[TBE.scala 114:59]
  wire [31:0] _GEN_884 = _T_111 ? _GEN_612 : _GEN_820; // @[TBE.scala 114:59]
  wire [31:0] _GEN_885 = _T_111 ? _GEN_613 : _GEN_821; // @[TBE.scala 114:59]
  wire [31:0] _GEN_886 = _T_111 ? _GEN_614 : _GEN_822; // @[TBE.scala 114:59]
  wire [31:0] _GEN_887 = _T_111 ? _GEN_615 : _GEN_823; // @[TBE.scala 114:59]
  wire [31:0] _GEN_888 = _T_111 ? _GEN_616 : _GEN_824; // @[TBE.scala 114:59]
  wire [31:0] _GEN_889 = _T_111 ? _GEN_617 : _GEN_825; // @[TBE.scala 114:59]
  wire [31:0] _GEN_890 = _T_111 ? _GEN_618 : _GEN_826; // @[TBE.scala 114:59]
  wire [31:0] _GEN_891 = _T_111 ? _GEN_619 : _GEN_827; // @[TBE.scala 114:59]
  wire [31:0] _GEN_892 = _T_111 ? _GEN_620 : _GEN_828; // @[TBE.scala 114:59]
  wire [31:0] _GEN_893 = _T_111 ? _GEN_621 : _GEN_829; // @[TBE.scala 114:59]
  wire [31:0] _GEN_894 = _T_111 ? _GEN_622 : _GEN_830; // @[TBE.scala 114:59]
  wire [31:0] _GEN_895 = _T_111 ? _GEN_623 : _GEN_831; // @[TBE.scala 114:59]
  wire [31:0] _GEN_896 = _T_111 ? _GEN_624 : _GEN_832; // @[TBE.scala 114:59]
  wire [31:0] _GEN_897 = _T_111 ? _GEN_625 : _GEN_833; // @[TBE.scala 114:59]
  wire [2:0] _GEN_898 = _T_111 ? _GEN_626 : _GEN_834; // @[TBE.scala 114:59]
  wire [2:0] _GEN_899 = _T_111 ? _GEN_627 : _GEN_835; // @[TBE.scala 114:59]
  wire [2:0] _GEN_900 = _T_111 ? _GEN_628 : _GEN_836; // @[TBE.scala 114:59]
  wire [2:0] _GEN_901 = _T_111 ? _GEN_629 : _GEN_837; // @[TBE.scala 114:59]
  wire [2:0] _GEN_902 = _T_111 ? _GEN_630 : _GEN_838; // @[TBE.scala 114:59]
  wire [2:0] _GEN_903 = _T_111 ? _GEN_631 : _GEN_839; // @[TBE.scala 114:59]
  wire [2:0] _GEN_904 = _T_111 ? _GEN_632 : _GEN_840; // @[TBE.scala 114:59]
  wire [2:0] _GEN_905 = _T_111 ? _GEN_633 : _GEN_841; // @[TBE.scala 114:59]
  wire [2:0] _GEN_906 = _T_111 ? _GEN_634 : _GEN_842; // @[TBE.scala 114:59]
  wire [2:0] _GEN_907 = _T_111 ? _GEN_635 : _GEN_843; // @[TBE.scala 114:59]
  wire [2:0] _GEN_908 = _T_111 ? _GEN_636 : _GEN_844; // @[TBE.scala 114:59]
  wire [2:0] _GEN_909 = _T_111 ? _GEN_637 : _GEN_845; // @[TBE.scala 114:59]
  wire [2:0] _GEN_910 = _T_111 ? _GEN_638 : _GEN_846; // @[TBE.scala 114:59]
  wire [2:0] _GEN_911 = _T_111 ? _GEN_639 : _GEN_847; // @[TBE.scala 114:59]
  wire [2:0] _GEN_912 = _T_111 ? _GEN_640 : _GEN_848; // @[TBE.scala 114:59]
  wire [2:0] _GEN_913 = _T_111 ? _GEN_641 : _GEN_849; // @[TBE.scala 114:59]
  wire [1:0] _GEN_914 = _T_111 ? _GEN_642 : _GEN_850; // @[TBE.scala 114:59]
  wire [1:0] _GEN_915 = _T_111 ? _GEN_643 : _GEN_851; // @[TBE.scala 114:59]
  wire [1:0] _GEN_916 = _T_111 ? _GEN_644 : _GEN_852; // @[TBE.scala 114:59]
  wire [1:0] _GEN_917 = _T_111 ? _GEN_645 : _GEN_853; // @[TBE.scala 114:59]
  wire [1:0] _GEN_918 = _T_111 ? _GEN_646 : _GEN_854; // @[TBE.scala 114:59]
  wire [1:0] _GEN_919 = _T_111 ? _GEN_647 : _GEN_855; // @[TBE.scala 114:59]
  wire [1:0] _GEN_920 = _T_111 ? _GEN_648 : _GEN_856; // @[TBE.scala 114:59]
  wire [1:0] _GEN_921 = _T_111 ? _GEN_649 : _GEN_857; // @[TBE.scala 114:59]
  wire [1:0] _GEN_922 = _T_111 ? _GEN_650 : _GEN_858; // @[TBE.scala 114:59]
  wire [1:0] _GEN_923 = _T_111 ? _GEN_651 : _GEN_859; // @[TBE.scala 114:59]
  wire [1:0] _GEN_924 = _T_111 ? _GEN_652 : _GEN_860; // @[TBE.scala 114:59]
  wire [1:0] _GEN_925 = _T_111 ? _GEN_653 : _GEN_861; // @[TBE.scala 114:59]
  wire [1:0] _GEN_926 = _T_111 ? _GEN_654 : _GEN_862; // @[TBE.scala 114:59]
  wire [1:0] _GEN_927 = _T_111 ? _GEN_655 : _GEN_863; // @[TBE.scala 114:59]
  wire [1:0] _GEN_928 = _T_111 ? _GEN_656 : _GEN_864; // @[TBE.scala 114:59]
  wire [1:0] _GEN_929 = _T_111 ? _GEN_657 : _GEN_865; // @[TBE.scala 114:59]
  wire [31:0] _GEN_930 = _T_111 ? _GEN_658 : _GEN_481; // @[TBE.scala 114:59]
  wire [31:0] _GEN_931 = _T_111 ? _GEN_659 : _GEN_482; // @[TBE.scala 114:59]
  wire [31:0] _GEN_932 = _T_111 ? _GEN_660 : _GEN_483; // @[TBE.scala 114:59]
  wire [31:0] _GEN_933 = _T_111 ? _GEN_661 : _GEN_484; // @[TBE.scala 114:59]
  wire [31:0] _GEN_934 = _T_111 ? _GEN_662 : _GEN_485; // @[TBE.scala 114:59]
  wire [31:0] _GEN_935 = _T_111 ? _GEN_663 : _GEN_486; // @[TBE.scala 114:59]
  wire [31:0] _GEN_936 = _T_111 ? _GEN_664 : _GEN_487; // @[TBE.scala 114:59]
  wire [31:0] _GEN_937 = _T_111 ? _GEN_665 : _GEN_488; // @[TBE.scala 114:59]
  wire [31:0] _GEN_938 = _T_111 ? _GEN_666 : _GEN_489; // @[TBE.scala 114:59]
  wire [31:0] _GEN_939 = _T_111 ? _GEN_667 : _GEN_490; // @[TBE.scala 114:59]
  wire [31:0] _GEN_940 = _T_111 ? _GEN_668 : _GEN_491; // @[TBE.scala 114:59]
  wire [31:0] _GEN_941 = _T_111 ? _GEN_669 : _GEN_492; // @[TBE.scala 114:59]
  wire [31:0] _GEN_942 = _T_111 ? _GEN_670 : _GEN_493; // @[TBE.scala 114:59]
  wire [31:0] _GEN_943 = _T_111 ? _GEN_671 : _GEN_494; // @[TBE.scala 114:59]
  wire [31:0] _GEN_944 = _T_111 ? _GEN_672 : _GEN_495; // @[TBE.scala 114:59]
  wire [31:0] _GEN_945 = _T_111 ? _GEN_673 : _GEN_496; // @[TBE.scala 114:59]
  wire  _T_269 = io_write_1_bits_command == 2'h1; // @[TBE.scala 136:44]
  wire  isAlloc_1 = _T_269 & io_write_1_valid; // @[TBE.scala 136:54]
  wire [31:0] _GEN_947 = isAlloc_1 ? _GEN_514 : _GEN_882; // @[TBE.scala 109:24]
  wire [31:0] _GEN_948 = isAlloc_1 ? _GEN_515 : _GEN_883; // @[TBE.scala 109:24]
  wire [31:0] _GEN_949 = isAlloc_1 ? _GEN_516 : _GEN_884; // @[TBE.scala 109:24]
  wire [31:0] _GEN_950 = isAlloc_1 ? _GEN_517 : _GEN_885; // @[TBE.scala 109:24]
  wire [31:0] _GEN_951 = isAlloc_1 ? _GEN_518 : _GEN_886; // @[TBE.scala 109:24]
  wire [31:0] _GEN_952 = isAlloc_1 ? _GEN_519 : _GEN_887; // @[TBE.scala 109:24]
  wire [31:0] _GEN_953 = isAlloc_1 ? _GEN_520 : _GEN_888; // @[TBE.scala 109:24]
  wire [31:0] _GEN_954 = isAlloc_1 ? _GEN_521 : _GEN_889; // @[TBE.scala 109:24]
  wire [31:0] _GEN_955 = isAlloc_1 ? _GEN_522 : _GEN_890; // @[TBE.scala 109:24]
  wire [31:0] _GEN_956 = isAlloc_1 ? _GEN_523 : _GEN_891; // @[TBE.scala 109:24]
  wire [31:0] _GEN_957 = isAlloc_1 ? _GEN_524 : _GEN_892; // @[TBE.scala 109:24]
  wire [31:0] _GEN_958 = isAlloc_1 ? _GEN_525 : _GEN_893; // @[TBE.scala 109:24]
  wire [31:0] _GEN_959 = isAlloc_1 ? _GEN_526 : _GEN_894; // @[TBE.scala 109:24]
  wire [31:0] _GEN_960 = isAlloc_1 ? _GEN_527 : _GEN_895; // @[TBE.scala 109:24]
  wire [31:0] _GEN_961 = isAlloc_1 ? _GEN_528 : _GEN_896; // @[TBE.scala 109:24]
  wire [31:0] _GEN_962 = isAlloc_1 ? _GEN_529 : _GEN_897; // @[TBE.scala 109:24]
  wire [2:0] _GEN_963 = isAlloc_1 ? _GEN_530 : _GEN_898; // @[TBE.scala 109:24]
  wire [2:0] _GEN_964 = isAlloc_1 ? _GEN_531 : _GEN_899; // @[TBE.scala 109:24]
  wire [2:0] _GEN_965 = isAlloc_1 ? _GEN_532 : _GEN_900; // @[TBE.scala 109:24]
  wire [2:0] _GEN_966 = isAlloc_1 ? _GEN_533 : _GEN_901; // @[TBE.scala 109:24]
  wire [2:0] _GEN_967 = isAlloc_1 ? _GEN_534 : _GEN_902; // @[TBE.scala 109:24]
  wire [2:0] _GEN_968 = isAlloc_1 ? _GEN_535 : _GEN_903; // @[TBE.scala 109:24]
  wire [2:0] _GEN_969 = isAlloc_1 ? _GEN_536 : _GEN_904; // @[TBE.scala 109:24]
  wire [2:0] _GEN_970 = isAlloc_1 ? _GEN_537 : _GEN_905; // @[TBE.scala 109:24]
  wire [2:0] _GEN_971 = isAlloc_1 ? _GEN_538 : _GEN_906; // @[TBE.scala 109:24]
  wire [2:0] _GEN_972 = isAlloc_1 ? _GEN_539 : _GEN_907; // @[TBE.scala 109:24]
  wire [2:0] _GEN_973 = isAlloc_1 ? _GEN_540 : _GEN_908; // @[TBE.scala 109:24]
  wire [2:0] _GEN_974 = isAlloc_1 ? _GEN_541 : _GEN_909; // @[TBE.scala 109:24]
  wire [2:0] _GEN_975 = isAlloc_1 ? _GEN_542 : _GEN_910; // @[TBE.scala 109:24]
  wire [2:0] _GEN_976 = isAlloc_1 ? _GEN_543 : _GEN_911; // @[TBE.scala 109:24]
  wire [2:0] _GEN_977 = isAlloc_1 ? _GEN_544 : _GEN_912; // @[TBE.scala 109:24]
  wire [2:0] _GEN_978 = isAlloc_1 ? _GEN_545 : _GEN_913; // @[TBE.scala 109:24]
  wire [1:0] _GEN_979 = isAlloc_1 ? _GEN_546 : _GEN_914; // @[TBE.scala 109:24]
  wire [1:0] _GEN_980 = isAlloc_1 ? _GEN_547 : _GEN_915; // @[TBE.scala 109:24]
  wire [1:0] _GEN_981 = isAlloc_1 ? _GEN_548 : _GEN_916; // @[TBE.scala 109:24]
  wire [1:0] _GEN_982 = isAlloc_1 ? _GEN_549 : _GEN_917; // @[TBE.scala 109:24]
  wire [1:0] _GEN_983 = isAlloc_1 ? _GEN_550 : _GEN_918; // @[TBE.scala 109:24]
  wire [1:0] _GEN_984 = isAlloc_1 ? _GEN_551 : _GEN_919; // @[TBE.scala 109:24]
  wire [1:0] _GEN_985 = isAlloc_1 ? _GEN_552 : _GEN_920; // @[TBE.scala 109:24]
  wire [1:0] _GEN_986 = isAlloc_1 ? _GEN_553 : _GEN_921; // @[TBE.scala 109:24]
  wire [1:0] _GEN_987 = isAlloc_1 ? _GEN_554 : _GEN_922; // @[TBE.scala 109:24]
  wire [1:0] _GEN_988 = isAlloc_1 ? _GEN_555 : _GEN_923; // @[TBE.scala 109:24]
  wire [1:0] _GEN_989 = isAlloc_1 ? _GEN_556 : _GEN_924; // @[TBE.scala 109:24]
  wire [1:0] _GEN_990 = isAlloc_1 ? _GEN_557 : _GEN_925; // @[TBE.scala 109:24]
  wire [1:0] _GEN_991 = isAlloc_1 ? _GEN_558 : _GEN_926; // @[TBE.scala 109:24]
  wire [1:0] _GEN_992 = isAlloc_1 ? _GEN_559 : _GEN_927; // @[TBE.scala 109:24]
  wire [1:0] _GEN_993 = isAlloc_1 ? _GEN_560 : _GEN_928; // @[TBE.scala 109:24]
  wire [1:0] _GEN_994 = isAlloc_1 ? _GEN_561 : _GEN_929; // @[TBE.scala 109:24]
  wire [31:0] _GEN_995 = isAlloc_1 ? _GEN_562 : _GEN_930; // @[TBE.scala 109:24]
  wire [31:0] _GEN_996 = isAlloc_1 ? _GEN_563 : _GEN_931; // @[TBE.scala 109:24]
  wire [31:0] _GEN_997 = isAlloc_1 ? _GEN_564 : _GEN_932; // @[TBE.scala 109:24]
  wire [31:0] _GEN_998 = isAlloc_1 ? _GEN_565 : _GEN_933; // @[TBE.scala 109:24]
  wire [31:0] _GEN_999 = isAlloc_1 ? _GEN_566 : _GEN_934; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1000 = isAlloc_1 ? _GEN_567 : _GEN_935; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1001 = isAlloc_1 ? _GEN_568 : _GEN_936; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1002 = isAlloc_1 ? _GEN_569 : _GEN_937; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1003 = isAlloc_1 ? _GEN_570 : _GEN_938; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1004 = isAlloc_1 ? _GEN_571 : _GEN_939; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1005 = isAlloc_1 ? _GEN_572 : _GEN_940; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1006 = isAlloc_1 ? _GEN_573 : _GEN_941; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1007 = isAlloc_1 ? _GEN_574 : _GEN_942; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1008 = isAlloc_1 ? _GEN_575 : _GEN_943; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1009 = isAlloc_1 ? _GEN_576 : _GEN_944; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1010 = isAlloc_1 ? _GEN_577 : _GEN_945; // @[TBE.scala 109:24]
  wire  _GEN_1011 = isAlloc_1 ? _GEN_578 : _GEN_866; // @[TBE.scala 109:24]
  wire  _GEN_1012 = isAlloc_1 ? _GEN_579 : _GEN_867; // @[TBE.scala 109:24]
  wire  _GEN_1013 = isAlloc_1 ? _GEN_580 : _GEN_868; // @[TBE.scala 109:24]
  wire  _GEN_1014 = isAlloc_1 ? _GEN_581 : _GEN_869; // @[TBE.scala 109:24]
  wire  _GEN_1015 = isAlloc_1 ? _GEN_582 : _GEN_870; // @[TBE.scala 109:24]
  wire  _GEN_1016 = isAlloc_1 ? _GEN_583 : _GEN_871; // @[TBE.scala 109:24]
  wire  _GEN_1017 = isAlloc_1 ? _GEN_584 : _GEN_872; // @[TBE.scala 109:24]
  wire  _GEN_1018 = isAlloc_1 ? _GEN_585 : _GEN_873; // @[TBE.scala 109:24]
  wire  _GEN_1019 = isAlloc_1 ? _GEN_586 : _GEN_874; // @[TBE.scala 109:24]
  wire  _GEN_1020 = isAlloc_1 ? _GEN_587 : _GEN_875; // @[TBE.scala 109:24]
  wire  _GEN_1021 = isAlloc_1 ? _GEN_588 : _GEN_876; // @[TBE.scala 109:24]
  wire  _GEN_1022 = isAlloc_1 ? _GEN_589 : _GEN_877; // @[TBE.scala 109:24]
  wire  _GEN_1023 = isAlloc_1 ? _GEN_590 : _GEN_878; // @[TBE.scala 109:24]
  wire  _GEN_1024 = isAlloc_1 ? _GEN_591 : _GEN_879; // @[TBE.scala 109:24]
  wire  _GEN_1025 = isAlloc_1 ? _GEN_592 : _GEN_880; // @[TBE.scala 109:24]
  wire  _GEN_1026 = isAlloc_1 ? _GEN_593 : _GEN_881; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1028 = 4'h0 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_947; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1029 = 4'h1 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_948; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1030 = 4'h2 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_949; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1031 = 4'h3 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_950; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1032 = 4'h4 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_951; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1033 = 4'h5 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_952; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1034 = 4'h6 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_953; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1035 = 4'h7 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_954; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1036 = 4'h8 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_955; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1037 = 4'h9 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_956; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1038 = 4'ha == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_957; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1039 = 4'hb == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_958; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1040 = 4'hc == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_959; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1041 = 4'hd == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_960; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1042 = 4'he == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_961; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1043 = 4'hf == idxAlloc[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_962; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1044 = 4'h0 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_963; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1045 = 4'h1 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_964; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1046 = 4'h2 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_965; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1047 = 4'h3 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_966; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1048 = 4'h4 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_967; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1049 = 4'h5 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_968; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1050 = 4'h6 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_969; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1051 = 4'h7 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_970; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1052 = 4'h8 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_971; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1053 = 4'h9 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_972; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1054 = 4'ha == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_973; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1055 = 4'hb == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_974; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1056 = 4'hc == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_975; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1057 = 4'hd == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_976; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1058 = 4'he == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_977; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1059 = 4'hf == idxAlloc[3:0] ? io_write_2_bits_inputTBE_way : _GEN_978; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1060 = 4'h0 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_979; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1061 = 4'h1 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_980; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1062 = 4'h2 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_981; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1063 = 4'h3 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_982; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1064 = 4'h4 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_983; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1065 = 4'h5 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_984; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1066 = 4'h6 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_985; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1067 = 4'h7 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_986; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1068 = 4'h8 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_987; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1069 = 4'h9 == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_988; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1070 = 4'ha == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_989; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1071 = 4'hb == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_990; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1072 = 4'hc == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_991; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1073 = 4'hd == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_992; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1074 = 4'he == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_993; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1075 = 4'hf == idxAlloc[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_994; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1076 = 4'h0 == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_995; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1077 = 4'h1 == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_996; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1078 = 4'h2 == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_997; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1079 = 4'h3 == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_998; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1080 = 4'h4 == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_999; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1081 = 4'h5 == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_1000; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1082 = 4'h6 == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_1001; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1083 = 4'h7 == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_1002; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1084 = 4'h8 == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_1003; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1085 = 4'h9 == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_1004; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1086 = 4'ha == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_1005; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1087 = 4'hb == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_1006; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1088 = 4'hc == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_1007; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1089 = 4'hd == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_1008; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1090 = 4'he == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_1009; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1091 = 4'hf == idxAlloc[3:0] ? io_write_2_bits_addr[31:0] : _GEN_1010; // @[TBE.scala 111:25]
  wire  _GEN_1092 = _GEN_4161 | _GEN_1011; // @[TBE.scala 112:26]
  wire  _GEN_1093 = _GEN_4162 | _GEN_1012; // @[TBE.scala 112:26]
  wire  _GEN_1094 = _GEN_4163 | _GEN_1013; // @[TBE.scala 112:26]
  wire  _GEN_1095 = _GEN_4164 | _GEN_1014; // @[TBE.scala 112:26]
  wire  _GEN_1096 = _GEN_4165 | _GEN_1015; // @[TBE.scala 112:26]
  wire  _GEN_1097 = _GEN_4166 | _GEN_1016; // @[TBE.scala 112:26]
  wire  _GEN_1098 = _GEN_4167 | _GEN_1017; // @[TBE.scala 112:26]
  wire  _GEN_1099 = _GEN_4168 | _GEN_1018; // @[TBE.scala 112:26]
  wire  _GEN_1100 = _GEN_4169 | _GEN_1019; // @[TBE.scala 112:26]
  wire  _GEN_1101 = _GEN_4170 | _GEN_1020; // @[TBE.scala 112:26]
  wire  _GEN_1102 = _GEN_4171 | _GEN_1021; // @[TBE.scala 112:26]
  wire  _GEN_1103 = _GEN_4172 | _GEN_1022; // @[TBE.scala 112:26]
  wire  _GEN_1104 = _GEN_4173 | _GEN_1023; // @[TBE.scala 112:26]
  wire  _GEN_1105 = _GEN_4174 | _GEN_1024; // @[TBE.scala 112:26]
  wire  _GEN_1106 = _GEN_4175 | _GEN_1025; // @[TBE.scala 112:26]
  wire  _GEN_1107 = _GEN_4176 | _GEN_1026; // @[TBE.scala 112:26]
  wire  _T_277 = io_write_2_bits_command == 2'h2; // @[TBE.scala 137:46]
  wire  isDealloc_2 = _T_277 & io_write_2_valid; // @[TBE.scala 137:58]
  wire  _T_133 = isDealloc_2 & finder_2_io_value_valid; // @[TBE.scala 114:31]
  wire [4:0] idxUpdate_2 = {{1'd0}, finder_2_io_value_bits}; // @[TBE.scala 73:23 TBE.scala 104:18]
  wire  _GEN_1108 = 4'h0 == idxUpdate_2[3:0] ? 1'h0 : _GEN_1011; // @[TBE.scala 115:30]
  wire  _GEN_1109 = 4'h1 == idxUpdate_2[3:0] ? 1'h0 : _GEN_1012; // @[TBE.scala 115:30]
  wire  _GEN_1110 = 4'h2 == idxUpdate_2[3:0] ? 1'h0 : _GEN_1013; // @[TBE.scala 115:30]
  wire  _GEN_1111 = 4'h3 == idxUpdate_2[3:0] ? 1'h0 : _GEN_1014; // @[TBE.scala 115:30]
  wire  _GEN_1112 = 4'h4 == idxUpdate_2[3:0] ? 1'h0 : _GEN_1015; // @[TBE.scala 115:30]
  wire  _GEN_1113 = 4'h5 == idxUpdate_2[3:0] ? 1'h0 : _GEN_1016; // @[TBE.scala 115:30]
  wire  _GEN_1114 = 4'h6 == idxUpdate_2[3:0] ? 1'h0 : _GEN_1017; // @[TBE.scala 115:30]
  wire  _GEN_1115 = 4'h7 == idxUpdate_2[3:0] ? 1'h0 : _GEN_1018; // @[TBE.scala 115:30]
  wire  _GEN_1116 = 4'h8 == idxUpdate_2[3:0] ? 1'h0 : _GEN_1019; // @[TBE.scala 115:30]
  wire  _GEN_1117 = 4'h9 == idxUpdate_2[3:0] ? 1'h0 : _GEN_1020; // @[TBE.scala 115:30]
  wire  _GEN_1118 = 4'ha == idxUpdate_2[3:0] ? 1'h0 : _GEN_1021; // @[TBE.scala 115:30]
  wire  _GEN_1119 = 4'hb == idxUpdate_2[3:0] ? 1'h0 : _GEN_1022; // @[TBE.scala 115:30]
  wire  _GEN_1120 = 4'hc == idxUpdate_2[3:0] ? 1'h0 : _GEN_1023; // @[TBE.scala 115:30]
  wire  _GEN_1121 = 4'hd == idxUpdate_2[3:0] ? 1'h0 : _GEN_1024; // @[TBE.scala 115:30]
  wire  _GEN_1122 = 4'he == idxUpdate_2[3:0] ? 1'h0 : _GEN_1025; // @[TBE.scala 115:30]
  wire  _GEN_1123 = 4'hf == idxUpdate_2[3:0] ? 1'h0 : _GEN_1026; // @[TBE.scala 115:30]
  wire [31:0] _GEN_1124 = 4'h0 == idxUpdate_2[3:0] ? 32'h0 : _GEN_947; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1125 = 4'h1 == idxUpdate_2[3:0] ? 32'h0 : _GEN_948; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1126 = 4'h2 == idxUpdate_2[3:0] ? 32'h0 : _GEN_949; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1127 = 4'h3 == idxUpdate_2[3:0] ? 32'h0 : _GEN_950; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1128 = 4'h4 == idxUpdate_2[3:0] ? 32'h0 : _GEN_951; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1129 = 4'h5 == idxUpdate_2[3:0] ? 32'h0 : _GEN_952; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1130 = 4'h6 == idxUpdate_2[3:0] ? 32'h0 : _GEN_953; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1131 = 4'h7 == idxUpdate_2[3:0] ? 32'h0 : _GEN_954; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1132 = 4'h8 == idxUpdate_2[3:0] ? 32'h0 : _GEN_955; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1133 = 4'h9 == idxUpdate_2[3:0] ? 32'h0 : _GEN_956; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1134 = 4'ha == idxUpdate_2[3:0] ? 32'h0 : _GEN_957; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1135 = 4'hb == idxUpdate_2[3:0] ? 32'h0 : _GEN_958; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1136 = 4'hc == idxUpdate_2[3:0] ? 32'h0 : _GEN_959; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1137 = 4'hd == idxUpdate_2[3:0] ? 32'h0 : _GEN_960; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1138 = 4'he == idxUpdate_2[3:0] ? 32'h0 : _GEN_961; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1139 = 4'hf == idxUpdate_2[3:0] ? 32'h0 : _GEN_962; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1140 = 4'h0 == idxUpdate_2[3:0] ? 3'h2 : _GEN_963; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1141 = 4'h1 == idxUpdate_2[3:0] ? 3'h2 : _GEN_964; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1142 = 4'h2 == idxUpdate_2[3:0] ? 3'h2 : _GEN_965; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1143 = 4'h3 == idxUpdate_2[3:0] ? 3'h2 : _GEN_966; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1144 = 4'h4 == idxUpdate_2[3:0] ? 3'h2 : _GEN_967; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1145 = 4'h5 == idxUpdate_2[3:0] ? 3'h2 : _GEN_968; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1146 = 4'h6 == idxUpdate_2[3:0] ? 3'h2 : _GEN_969; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1147 = 4'h7 == idxUpdate_2[3:0] ? 3'h2 : _GEN_970; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1148 = 4'h8 == idxUpdate_2[3:0] ? 3'h2 : _GEN_971; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1149 = 4'h9 == idxUpdate_2[3:0] ? 3'h2 : _GEN_972; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1150 = 4'ha == idxUpdate_2[3:0] ? 3'h2 : _GEN_973; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1151 = 4'hb == idxUpdate_2[3:0] ? 3'h2 : _GEN_974; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1152 = 4'hc == idxUpdate_2[3:0] ? 3'h2 : _GEN_975; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1153 = 4'hd == idxUpdate_2[3:0] ? 3'h2 : _GEN_976; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1154 = 4'he == idxUpdate_2[3:0] ? 3'h2 : _GEN_977; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1155 = 4'hf == idxUpdate_2[3:0] ? 3'h2 : _GEN_978; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1156 = 4'h0 == idxUpdate_2[3:0] ? 2'h0 : _GEN_979; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1157 = 4'h1 == idxUpdate_2[3:0] ? 2'h0 : _GEN_980; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1158 = 4'h2 == idxUpdate_2[3:0] ? 2'h0 : _GEN_981; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1159 = 4'h3 == idxUpdate_2[3:0] ? 2'h0 : _GEN_982; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1160 = 4'h4 == idxUpdate_2[3:0] ? 2'h0 : _GEN_983; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1161 = 4'h5 == idxUpdate_2[3:0] ? 2'h0 : _GEN_984; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1162 = 4'h6 == idxUpdate_2[3:0] ? 2'h0 : _GEN_985; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1163 = 4'h7 == idxUpdate_2[3:0] ? 2'h0 : _GEN_986; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1164 = 4'h8 == idxUpdate_2[3:0] ? 2'h0 : _GEN_987; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1165 = 4'h9 == idxUpdate_2[3:0] ? 2'h0 : _GEN_988; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1166 = 4'ha == idxUpdate_2[3:0] ? 2'h0 : _GEN_989; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1167 = 4'hb == idxUpdate_2[3:0] ? 2'h0 : _GEN_990; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1168 = 4'hc == idxUpdate_2[3:0] ? 2'h0 : _GEN_991; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1169 = 4'hd == idxUpdate_2[3:0] ? 2'h0 : _GEN_992; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1170 = 4'he == idxUpdate_2[3:0] ? 2'h0 : _GEN_993; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1171 = 4'hf == idxUpdate_2[3:0] ? 2'h0 : _GEN_994; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1172 = 4'h0 == idxUpdate_2[3:0] ? 32'h0 : _GEN_995; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1173 = 4'h1 == idxUpdate_2[3:0] ? 32'h0 : _GEN_996; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1174 = 4'h2 == idxUpdate_2[3:0] ? 32'h0 : _GEN_997; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1175 = 4'h3 == idxUpdate_2[3:0] ? 32'h0 : _GEN_998; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1176 = 4'h4 == idxUpdate_2[3:0] ? 32'h0 : _GEN_999; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1177 = 4'h5 == idxUpdate_2[3:0] ? 32'h0 : _GEN_1000; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1178 = 4'h6 == idxUpdate_2[3:0] ? 32'h0 : _GEN_1001; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1179 = 4'h7 == idxUpdate_2[3:0] ? 32'h0 : _GEN_1002; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1180 = 4'h8 == idxUpdate_2[3:0] ? 32'h0 : _GEN_1003; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1181 = 4'h9 == idxUpdate_2[3:0] ? 32'h0 : _GEN_1004; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1182 = 4'ha == idxUpdate_2[3:0] ? 32'h0 : _GEN_1005; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1183 = 4'hb == idxUpdate_2[3:0] ? 32'h0 : _GEN_1006; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1184 = 4'hc == idxUpdate_2[3:0] ? 32'h0 : _GEN_1007; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1185 = 4'hd == idxUpdate_2[3:0] ? 32'h0 : _GEN_1008; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1186 = 4'he == idxUpdate_2[3:0] ? 32'h0 : _GEN_1009; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1187 = 4'hf == idxUpdate_2[3:0] ? 32'h0 : _GEN_1010; // @[TBE.scala 117:29]
  wire  _T_279 = io_write_2_bits_command == 2'h3; // @[TBE.scala 138:44]
  wire  isWrite_2 = _T_279 & io_write_2_valid; // @[TBE.scala 138:55]
  wire  _T_141 = isWrite_2 & finder_2_io_value_valid; // @[TBE.scala 119:29]
  wire  _T_142 = ~io_write_2_bits_mask; // @[TBE.scala 120:35]
  wire [31:0] _GEN_1188 = 4'h0 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_947; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1189 = 4'h1 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_948; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1190 = 4'h2 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_949; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1191 = 4'h3 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_950; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1192 = 4'h4 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_951; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1193 = 4'h5 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_952; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1194 = 4'h6 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_953; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1195 = 4'h7 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_954; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1196 = 4'h8 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_955; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1197 = 4'h9 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_956; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1198 = 4'ha == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_957; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1199 = 4'hb == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_958; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1200 = 4'hc == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_959; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1201 = 4'hd == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_960; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1202 = 4'he == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_961; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1203 = 4'hf == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_fields_0 : _GEN_962; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1209 = 4'h1 == idxUpdate_2[3:0] ? TBEMemory_1_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1212 = 4'h2 == idxUpdate_2[3:0] ? TBEMemory_2_fields_0 : _GEN_1209; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1215 = 4'h3 == idxUpdate_2[3:0] ? TBEMemory_3_fields_0 : _GEN_1212; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1218 = 4'h4 == idxUpdate_2[3:0] ? TBEMemory_4_fields_0 : _GEN_1215; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1221 = 4'h5 == idxUpdate_2[3:0] ? TBEMemory_5_fields_0 : _GEN_1218; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1224 = 4'h6 == idxUpdate_2[3:0] ? TBEMemory_6_fields_0 : _GEN_1221; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1227 = 4'h7 == idxUpdate_2[3:0] ? TBEMemory_7_fields_0 : _GEN_1224; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1230 = 4'h8 == idxUpdate_2[3:0] ? TBEMemory_8_fields_0 : _GEN_1227; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1233 = 4'h9 == idxUpdate_2[3:0] ? TBEMemory_9_fields_0 : _GEN_1230; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1236 = 4'ha == idxUpdate_2[3:0] ? TBEMemory_10_fields_0 : _GEN_1233; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1239 = 4'hb == idxUpdate_2[3:0] ? TBEMemory_11_fields_0 : _GEN_1236; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1242 = 4'hc == idxUpdate_2[3:0] ? TBEMemory_12_fields_0 : _GEN_1239; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1245 = 4'hd == idxUpdate_2[3:0] ? TBEMemory_13_fields_0 : _GEN_1242; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1248 = 4'he == idxUpdate_2[3:0] ? TBEMemory_14_fields_0 : _GEN_1245; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1251 = 4'hf == idxUpdate_2[3:0] ? TBEMemory_15_fields_0 : _GEN_1248; // @[TBE.scala 122:15]
  wire [2:0] _GEN_1252 = 4'h0 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_963; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1253 = 4'h1 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_964; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1254 = 4'h2 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_965; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1255 = 4'h3 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_966; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1256 = 4'h4 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_967; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1257 = 4'h5 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_968; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1258 = 4'h6 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_969; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1259 = 4'h7 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_970; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1260 = 4'h8 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_971; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1261 = 4'h9 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_972; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1262 = 4'ha == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_973; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1263 = 4'hb == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_974; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1264 = 4'hc == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_975; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1265 = 4'hd == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_976; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1266 = 4'he == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_977; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1267 = 4'hf == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_way : _GEN_978; // @[TBE.scala 124:37]
  wire [1:0] _GEN_1268 = 4'h0 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_979; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1269 = 4'h1 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_980; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1270 = 4'h2 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_981; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1271 = 4'h3 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_982; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1272 = 4'h4 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_983; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1273 = 4'h5 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_984; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1274 = 4'h6 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_985; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1275 = 4'h7 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_986; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1276 = 4'h8 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_987; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1277 = 4'h9 == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_988; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1278 = 4'ha == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_989; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1279 = 4'hb == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_990; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1280 = 4'hc == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_991; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1281 = 4'hd == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_992; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1282 = 4'he == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_993; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1283 = 4'hf == idxUpdate_2[3:0] ? io_write_2_bits_inputTBE_state_state : _GEN_994; // @[TBE.scala 125:39]
  wire [31:0] _GEN_1284 = _T_142 ? _GEN_1188 : _GEN_947; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1285 = _T_142 ? _GEN_1189 : _GEN_948; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1286 = _T_142 ? _GEN_1190 : _GEN_949; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1287 = _T_142 ? _GEN_1191 : _GEN_950; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1288 = _T_142 ? _GEN_1192 : _GEN_951; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1289 = _T_142 ? _GEN_1193 : _GEN_952; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1290 = _T_142 ? _GEN_1194 : _GEN_953; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1291 = _T_142 ? _GEN_1195 : _GEN_954; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1292 = _T_142 ? _GEN_1196 : _GEN_955; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1293 = _T_142 ? _GEN_1197 : _GEN_956; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1294 = _T_142 ? _GEN_1198 : _GEN_957; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1295 = _T_142 ? _GEN_1199 : _GEN_958; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1296 = _T_142 ? _GEN_1200 : _GEN_959; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1297 = _T_142 ? _GEN_1201 : _GEN_960; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1298 = _T_142 ? _GEN_1202 : _GEN_961; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1299 = _T_142 ? _GEN_1203 : _GEN_962; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1300 = _T_142 ? _GEN_963 : _GEN_1252; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1301 = _T_142 ? _GEN_964 : _GEN_1253; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1302 = _T_142 ? _GEN_965 : _GEN_1254; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1303 = _T_142 ? _GEN_966 : _GEN_1255; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1304 = _T_142 ? _GEN_967 : _GEN_1256; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1305 = _T_142 ? _GEN_968 : _GEN_1257; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1306 = _T_142 ? _GEN_969 : _GEN_1258; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1307 = _T_142 ? _GEN_970 : _GEN_1259; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1308 = _T_142 ? _GEN_971 : _GEN_1260; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1309 = _T_142 ? _GEN_972 : _GEN_1261; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1310 = _T_142 ? _GEN_973 : _GEN_1262; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1311 = _T_142 ? _GEN_974 : _GEN_1263; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1312 = _T_142 ? _GEN_975 : _GEN_1264; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1313 = _T_142 ? _GEN_976 : _GEN_1265; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1314 = _T_142 ? _GEN_977 : _GEN_1266; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1315 = _T_142 ? _GEN_978 : _GEN_1267; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1316 = _T_142 ? _GEN_979 : _GEN_1268; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1317 = _T_142 ? _GEN_980 : _GEN_1269; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1318 = _T_142 ? _GEN_981 : _GEN_1270; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1319 = _T_142 ? _GEN_982 : _GEN_1271; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1320 = _T_142 ? _GEN_983 : _GEN_1272; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1321 = _T_142 ? _GEN_984 : _GEN_1273; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1322 = _T_142 ? _GEN_985 : _GEN_1274; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1323 = _T_142 ? _GEN_986 : _GEN_1275; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1324 = _T_142 ? _GEN_987 : _GEN_1276; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1325 = _T_142 ? _GEN_988 : _GEN_1277; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1326 = _T_142 ? _GEN_989 : _GEN_1278; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1327 = _T_142 ? _GEN_990 : _GEN_1279; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1328 = _T_142 ? _GEN_991 : _GEN_1280; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1329 = _T_142 ? _GEN_992 : _GEN_1281; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1330 = _T_142 ? _GEN_993 : _GEN_1282; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1331 = _T_142 ? _GEN_994 : _GEN_1283; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1332 = _T_141 ? _GEN_1284 : _GEN_947; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1333 = _T_141 ? _GEN_1285 : _GEN_948; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1334 = _T_141 ? _GEN_1286 : _GEN_949; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1335 = _T_141 ? _GEN_1287 : _GEN_950; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1336 = _T_141 ? _GEN_1288 : _GEN_951; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1337 = _T_141 ? _GEN_1289 : _GEN_952; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1338 = _T_141 ? _GEN_1290 : _GEN_953; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1339 = _T_141 ? _GEN_1291 : _GEN_954; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1340 = _T_141 ? _GEN_1292 : _GEN_955; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1341 = _T_141 ? _GEN_1293 : _GEN_956; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1342 = _T_141 ? _GEN_1294 : _GEN_957; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1343 = _T_141 ? _GEN_1295 : _GEN_958; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1344 = _T_141 ? _GEN_1296 : _GEN_959; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1345 = _T_141 ? _GEN_1297 : _GEN_960; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1346 = _T_141 ? _GEN_1298 : _GEN_961; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1347 = _T_141 ? _GEN_1299 : _GEN_962; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1348 = _T_141 ? _GEN_1300 : _GEN_963; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1349 = _T_141 ? _GEN_1301 : _GEN_964; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1350 = _T_141 ? _GEN_1302 : _GEN_965; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1351 = _T_141 ? _GEN_1303 : _GEN_966; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1352 = _T_141 ? _GEN_1304 : _GEN_967; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1353 = _T_141 ? _GEN_1305 : _GEN_968; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1354 = _T_141 ? _GEN_1306 : _GEN_969; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1355 = _T_141 ? _GEN_1307 : _GEN_970; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1356 = _T_141 ? _GEN_1308 : _GEN_971; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1357 = _T_141 ? _GEN_1309 : _GEN_972; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1358 = _T_141 ? _GEN_1310 : _GEN_973; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1359 = _T_141 ? _GEN_1311 : _GEN_974; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1360 = _T_141 ? _GEN_1312 : _GEN_975; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1361 = _T_141 ? _GEN_1313 : _GEN_976; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1362 = _T_141 ? _GEN_1314 : _GEN_977; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1363 = _T_141 ? _GEN_1315 : _GEN_978; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1364 = _T_141 ? _GEN_1316 : _GEN_979; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1365 = _T_141 ? _GEN_1317 : _GEN_980; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1366 = _T_141 ? _GEN_1318 : _GEN_981; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1367 = _T_141 ? _GEN_1319 : _GEN_982; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1368 = _T_141 ? _GEN_1320 : _GEN_983; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1369 = _T_141 ? _GEN_1321 : _GEN_984; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1370 = _T_141 ? _GEN_1322 : _GEN_985; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1371 = _T_141 ? _GEN_1323 : _GEN_986; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1372 = _T_141 ? _GEN_1324 : _GEN_987; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1373 = _T_141 ? _GEN_1325 : _GEN_988; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1374 = _T_141 ? _GEN_1326 : _GEN_989; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1375 = _T_141 ? _GEN_1327 : _GEN_990; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1376 = _T_141 ? _GEN_1328 : _GEN_991; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1377 = _T_141 ? _GEN_1329 : _GEN_992; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1378 = _T_141 ? _GEN_1330 : _GEN_993; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1379 = _T_141 ? _GEN_1331 : _GEN_994; // @[TBE.scala 119:57]
  wire  _GEN_1380 = _T_133 ? _GEN_1108 : _GEN_1011; // @[TBE.scala 114:59]
  wire  _GEN_1381 = _T_133 ? _GEN_1109 : _GEN_1012; // @[TBE.scala 114:59]
  wire  _GEN_1382 = _T_133 ? _GEN_1110 : _GEN_1013; // @[TBE.scala 114:59]
  wire  _GEN_1383 = _T_133 ? _GEN_1111 : _GEN_1014; // @[TBE.scala 114:59]
  wire  _GEN_1384 = _T_133 ? _GEN_1112 : _GEN_1015; // @[TBE.scala 114:59]
  wire  _GEN_1385 = _T_133 ? _GEN_1113 : _GEN_1016; // @[TBE.scala 114:59]
  wire  _GEN_1386 = _T_133 ? _GEN_1114 : _GEN_1017; // @[TBE.scala 114:59]
  wire  _GEN_1387 = _T_133 ? _GEN_1115 : _GEN_1018; // @[TBE.scala 114:59]
  wire  _GEN_1388 = _T_133 ? _GEN_1116 : _GEN_1019; // @[TBE.scala 114:59]
  wire  _GEN_1389 = _T_133 ? _GEN_1117 : _GEN_1020; // @[TBE.scala 114:59]
  wire  _GEN_1390 = _T_133 ? _GEN_1118 : _GEN_1021; // @[TBE.scala 114:59]
  wire  _GEN_1391 = _T_133 ? _GEN_1119 : _GEN_1022; // @[TBE.scala 114:59]
  wire  _GEN_1392 = _T_133 ? _GEN_1120 : _GEN_1023; // @[TBE.scala 114:59]
  wire  _GEN_1393 = _T_133 ? _GEN_1121 : _GEN_1024; // @[TBE.scala 114:59]
  wire  _GEN_1394 = _T_133 ? _GEN_1122 : _GEN_1025; // @[TBE.scala 114:59]
  wire  _GEN_1395 = _T_133 ? _GEN_1123 : _GEN_1026; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1396 = _T_133 ? _GEN_1124 : _GEN_1332; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1397 = _T_133 ? _GEN_1125 : _GEN_1333; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1398 = _T_133 ? _GEN_1126 : _GEN_1334; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1399 = _T_133 ? _GEN_1127 : _GEN_1335; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1400 = _T_133 ? _GEN_1128 : _GEN_1336; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1401 = _T_133 ? _GEN_1129 : _GEN_1337; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1402 = _T_133 ? _GEN_1130 : _GEN_1338; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1403 = _T_133 ? _GEN_1131 : _GEN_1339; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1404 = _T_133 ? _GEN_1132 : _GEN_1340; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1405 = _T_133 ? _GEN_1133 : _GEN_1341; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1406 = _T_133 ? _GEN_1134 : _GEN_1342; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1407 = _T_133 ? _GEN_1135 : _GEN_1343; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1408 = _T_133 ? _GEN_1136 : _GEN_1344; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1409 = _T_133 ? _GEN_1137 : _GEN_1345; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1410 = _T_133 ? _GEN_1138 : _GEN_1346; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1411 = _T_133 ? _GEN_1139 : _GEN_1347; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1412 = _T_133 ? _GEN_1140 : _GEN_1348; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1413 = _T_133 ? _GEN_1141 : _GEN_1349; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1414 = _T_133 ? _GEN_1142 : _GEN_1350; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1415 = _T_133 ? _GEN_1143 : _GEN_1351; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1416 = _T_133 ? _GEN_1144 : _GEN_1352; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1417 = _T_133 ? _GEN_1145 : _GEN_1353; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1418 = _T_133 ? _GEN_1146 : _GEN_1354; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1419 = _T_133 ? _GEN_1147 : _GEN_1355; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1420 = _T_133 ? _GEN_1148 : _GEN_1356; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1421 = _T_133 ? _GEN_1149 : _GEN_1357; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1422 = _T_133 ? _GEN_1150 : _GEN_1358; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1423 = _T_133 ? _GEN_1151 : _GEN_1359; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1424 = _T_133 ? _GEN_1152 : _GEN_1360; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1425 = _T_133 ? _GEN_1153 : _GEN_1361; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1426 = _T_133 ? _GEN_1154 : _GEN_1362; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1427 = _T_133 ? _GEN_1155 : _GEN_1363; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1428 = _T_133 ? _GEN_1156 : _GEN_1364; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1429 = _T_133 ? _GEN_1157 : _GEN_1365; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1430 = _T_133 ? _GEN_1158 : _GEN_1366; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1431 = _T_133 ? _GEN_1159 : _GEN_1367; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1432 = _T_133 ? _GEN_1160 : _GEN_1368; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1433 = _T_133 ? _GEN_1161 : _GEN_1369; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1434 = _T_133 ? _GEN_1162 : _GEN_1370; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1435 = _T_133 ? _GEN_1163 : _GEN_1371; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1436 = _T_133 ? _GEN_1164 : _GEN_1372; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1437 = _T_133 ? _GEN_1165 : _GEN_1373; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1438 = _T_133 ? _GEN_1166 : _GEN_1374; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1439 = _T_133 ? _GEN_1167 : _GEN_1375; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1440 = _T_133 ? _GEN_1168 : _GEN_1376; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1441 = _T_133 ? _GEN_1169 : _GEN_1377; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1442 = _T_133 ? _GEN_1170 : _GEN_1378; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1443 = _T_133 ? _GEN_1171 : _GEN_1379; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1444 = _T_133 ? _GEN_1172 : _GEN_995; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1445 = _T_133 ? _GEN_1173 : _GEN_996; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1446 = _T_133 ? _GEN_1174 : _GEN_997; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1447 = _T_133 ? _GEN_1175 : _GEN_998; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1448 = _T_133 ? _GEN_1176 : _GEN_999; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1449 = _T_133 ? _GEN_1177 : _GEN_1000; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1450 = _T_133 ? _GEN_1178 : _GEN_1001; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1451 = _T_133 ? _GEN_1179 : _GEN_1002; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1452 = _T_133 ? _GEN_1180 : _GEN_1003; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1453 = _T_133 ? _GEN_1181 : _GEN_1004; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1454 = _T_133 ? _GEN_1182 : _GEN_1005; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1455 = _T_133 ? _GEN_1183 : _GEN_1006; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1456 = _T_133 ? _GEN_1184 : _GEN_1007; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1457 = _T_133 ? _GEN_1185 : _GEN_1008; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1458 = _T_133 ? _GEN_1186 : _GEN_1009; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1459 = _T_133 ? _GEN_1187 : _GEN_1010; // @[TBE.scala 114:59]
  wire  _T_275 = io_write_2_bits_command == 2'h1; // @[TBE.scala 136:44]
  wire  isAlloc_2 = _T_275 & io_write_2_valid; // @[TBE.scala 136:54]
  wire [31:0] _GEN_1461 = isAlloc_2 ? _GEN_1028 : _GEN_1396; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1462 = isAlloc_2 ? _GEN_1029 : _GEN_1397; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1463 = isAlloc_2 ? _GEN_1030 : _GEN_1398; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1464 = isAlloc_2 ? _GEN_1031 : _GEN_1399; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1465 = isAlloc_2 ? _GEN_1032 : _GEN_1400; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1466 = isAlloc_2 ? _GEN_1033 : _GEN_1401; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1467 = isAlloc_2 ? _GEN_1034 : _GEN_1402; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1468 = isAlloc_2 ? _GEN_1035 : _GEN_1403; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1469 = isAlloc_2 ? _GEN_1036 : _GEN_1404; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1470 = isAlloc_2 ? _GEN_1037 : _GEN_1405; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1471 = isAlloc_2 ? _GEN_1038 : _GEN_1406; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1472 = isAlloc_2 ? _GEN_1039 : _GEN_1407; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1473 = isAlloc_2 ? _GEN_1040 : _GEN_1408; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1474 = isAlloc_2 ? _GEN_1041 : _GEN_1409; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1475 = isAlloc_2 ? _GEN_1042 : _GEN_1410; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1476 = isAlloc_2 ? _GEN_1043 : _GEN_1411; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1477 = isAlloc_2 ? _GEN_1044 : _GEN_1412; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1478 = isAlloc_2 ? _GEN_1045 : _GEN_1413; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1479 = isAlloc_2 ? _GEN_1046 : _GEN_1414; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1480 = isAlloc_2 ? _GEN_1047 : _GEN_1415; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1481 = isAlloc_2 ? _GEN_1048 : _GEN_1416; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1482 = isAlloc_2 ? _GEN_1049 : _GEN_1417; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1483 = isAlloc_2 ? _GEN_1050 : _GEN_1418; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1484 = isAlloc_2 ? _GEN_1051 : _GEN_1419; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1485 = isAlloc_2 ? _GEN_1052 : _GEN_1420; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1486 = isAlloc_2 ? _GEN_1053 : _GEN_1421; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1487 = isAlloc_2 ? _GEN_1054 : _GEN_1422; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1488 = isAlloc_2 ? _GEN_1055 : _GEN_1423; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1489 = isAlloc_2 ? _GEN_1056 : _GEN_1424; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1490 = isAlloc_2 ? _GEN_1057 : _GEN_1425; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1491 = isAlloc_2 ? _GEN_1058 : _GEN_1426; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1492 = isAlloc_2 ? _GEN_1059 : _GEN_1427; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1493 = isAlloc_2 ? _GEN_1060 : _GEN_1428; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1494 = isAlloc_2 ? _GEN_1061 : _GEN_1429; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1495 = isAlloc_2 ? _GEN_1062 : _GEN_1430; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1496 = isAlloc_2 ? _GEN_1063 : _GEN_1431; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1497 = isAlloc_2 ? _GEN_1064 : _GEN_1432; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1498 = isAlloc_2 ? _GEN_1065 : _GEN_1433; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1499 = isAlloc_2 ? _GEN_1066 : _GEN_1434; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1500 = isAlloc_2 ? _GEN_1067 : _GEN_1435; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1501 = isAlloc_2 ? _GEN_1068 : _GEN_1436; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1502 = isAlloc_2 ? _GEN_1069 : _GEN_1437; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1503 = isAlloc_2 ? _GEN_1070 : _GEN_1438; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1504 = isAlloc_2 ? _GEN_1071 : _GEN_1439; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1505 = isAlloc_2 ? _GEN_1072 : _GEN_1440; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1506 = isAlloc_2 ? _GEN_1073 : _GEN_1441; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1507 = isAlloc_2 ? _GEN_1074 : _GEN_1442; // @[TBE.scala 109:24]
  wire [1:0] _GEN_1508 = isAlloc_2 ? _GEN_1075 : _GEN_1443; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1509 = isAlloc_2 ? _GEN_1076 : _GEN_1444; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1510 = isAlloc_2 ? _GEN_1077 : _GEN_1445; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1511 = isAlloc_2 ? _GEN_1078 : _GEN_1446; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1512 = isAlloc_2 ? _GEN_1079 : _GEN_1447; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1513 = isAlloc_2 ? _GEN_1080 : _GEN_1448; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1514 = isAlloc_2 ? _GEN_1081 : _GEN_1449; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1515 = isAlloc_2 ? _GEN_1082 : _GEN_1450; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1516 = isAlloc_2 ? _GEN_1083 : _GEN_1451; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1517 = isAlloc_2 ? _GEN_1084 : _GEN_1452; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1518 = isAlloc_2 ? _GEN_1085 : _GEN_1453; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1519 = isAlloc_2 ? _GEN_1086 : _GEN_1454; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1520 = isAlloc_2 ? _GEN_1087 : _GEN_1455; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1521 = isAlloc_2 ? _GEN_1088 : _GEN_1456; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1522 = isAlloc_2 ? _GEN_1089 : _GEN_1457; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1523 = isAlloc_2 ? _GEN_1090 : _GEN_1458; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1524 = isAlloc_2 ? _GEN_1091 : _GEN_1459; // @[TBE.scala 109:24]
  wire  _GEN_1525 = isAlloc_2 ? _GEN_1092 : _GEN_1380; // @[TBE.scala 109:24]
  wire  _GEN_1526 = isAlloc_2 ? _GEN_1093 : _GEN_1381; // @[TBE.scala 109:24]
  wire  _GEN_1527 = isAlloc_2 ? _GEN_1094 : _GEN_1382; // @[TBE.scala 109:24]
  wire  _GEN_1528 = isAlloc_2 ? _GEN_1095 : _GEN_1383; // @[TBE.scala 109:24]
  wire  _GEN_1529 = isAlloc_2 ? _GEN_1096 : _GEN_1384; // @[TBE.scala 109:24]
  wire  _GEN_1530 = isAlloc_2 ? _GEN_1097 : _GEN_1385; // @[TBE.scala 109:24]
  wire  _GEN_1531 = isAlloc_2 ? _GEN_1098 : _GEN_1386; // @[TBE.scala 109:24]
  wire  _GEN_1532 = isAlloc_2 ? _GEN_1099 : _GEN_1387; // @[TBE.scala 109:24]
  wire  _GEN_1533 = isAlloc_2 ? _GEN_1100 : _GEN_1388; // @[TBE.scala 109:24]
  wire  _GEN_1534 = isAlloc_2 ? _GEN_1101 : _GEN_1389; // @[TBE.scala 109:24]
  wire  _GEN_1535 = isAlloc_2 ? _GEN_1102 : _GEN_1390; // @[TBE.scala 109:24]
  wire  _GEN_1536 = isAlloc_2 ? _GEN_1103 : _GEN_1391; // @[TBE.scala 109:24]
  wire  _GEN_1537 = isAlloc_2 ? _GEN_1104 : _GEN_1392; // @[TBE.scala 109:24]
  wire  _GEN_1538 = isAlloc_2 ? _GEN_1105 : _GEN_1393; // @[TBE.scala 109:24]
  wire  _GEN_1539 = isAlloc_2 ? _GEN_1106 : _GEN_1394; // @[TBE.scala 109:24]
  wire  _GEN_1540 = isAlloc_2 ? _GEN_1107 : _GEN_1395; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1542 = 4'h0 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1461; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1543 = 4'h1 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1462; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1544 = 4'h2 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1463; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1545 = 4'h3 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1464; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1546 = 4'h4 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1465; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1547 = 4'h5 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1466; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1548 = 4'h6 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1467; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1549 = 4'h7 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1468; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1550 = 4'h8 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1469; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1551 = 4'h9 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1470; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1552 = 4'ha == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1471; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1553 = 4'hb == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1472; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1554 = 4'hc == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1473; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1555 = 4'hd == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1474; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1556 = 4'he == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1475; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1557 = 4'hf == idxAlloc[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1476; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1558 = 4'h0 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1477; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1559 = 4'h1 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1478; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1560 = 4'h2 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1479; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1561 = 4'h3 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1480; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1562 = 4'h4 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1481; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1563 = 4'h5 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1482; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1564 = 4'h6 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1483; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1565 = 4'h7 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1484; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1566 = 4'h8 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1485; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1567 = 4'h9 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1486; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1568 = 4'ha == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1487; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1569 = 4'hb == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1488; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1570 = 4'hc == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1489; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1571 = 4'hd == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1490; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1572 = 4'he == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1491; // @[TBE.scala 110:27]
  wire [2:0] _GEN_1573 = 4'hf == idxAlloc[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1492; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1574 = 4'h0 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1493; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1575 = 4'h1 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1494; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1576 = 4'h2 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1495; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1577 = 4'h3 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1496; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1578 = 4'h4 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1497; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1579 = 4'h5 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1498; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1580 = 4'h6 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1499; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1581 = 4'h7 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1500; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1582 = 4'h8 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1501; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1583 = 4'h9 == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1502; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1584 = 4'ha == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1503; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1585 = 4'hb == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1504; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1586 = 4'hc == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1505; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1587 = 4'hd == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1506; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1588 = 4'he == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1507; // @[TBE.scala 110:27]
  wire [1:0] _GEN_1589 = 4'hf == idxAlloc[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1508; // @[TBE.scala 110:27]
  wire [31:0] _GEN_1590 = 4'h0 == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1509; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1591 = 4'h1 == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1510; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1592 = 4'h2 == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1511; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1593 = 4'h3 == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1512; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1594 = 4'h4 == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1513; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1595 = 4'h5 == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1514; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1596 = 4'h6 == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1515; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1597 = 4'h7 == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1516; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1598 = 4'h8 == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1517; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1599 = 4'h9 == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1518; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1600 = 4'ha == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1519; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1601 = 4'hb == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1520; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1602 = 4'hc == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1521; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1603 = 4'hd == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1522; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1604 = 4'he == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1523; // @[TBE.scala 111:25]
  wire [31:0] _GEN_1605 = 4'hf == idxAlloc[3:0] ? io_write_3_bits_addr[31:0] : _GEN_1524; // @[TBE.scala 111:25]
  wire  _GEN_1606 = _GEN_4161 | _GEN_1525; // @[TBE.scala 112:26]
  wire  _GEN_1607 = _GEN_4162 | _GEN_1526; // @[TBE.scala 112:26]
  wire  _GEN_1608 = _GEN_4163 | _GEN_1527; // @[TBE.scala 112:26]
  wire  _GEN_1609 = _GEN_4164 | _GEN_1528; // @[TBE.scala 112:26]
  wire  _GEN_1610 = _GEN_4165 | _GEN_1529; // @[TBE.scala 112:26]
  wire  _GEN_1611 = _GEN_4166 | _GEN_1530; // @[TBE.scala 112:26]
  wire  _GEN_1612 = _GEN_4167 | _GEN_1531; // @[TBE.scala 112:26]
  wire  _GEN_1613 = _GEN_4168 | _GEN_1532; // @[TBE.scala 112:26]
  wire  _GEN_1614 = _GEN_4169 | _GEN_1533; // @[TBE.scala 112:26]
  wire  _GEN_1615 = _GEN_4170 | _GEN_1534; // @[TBE.scala 112:26]
  wire  _GEN_1616 = _GEN_4171 | _GEN_1535; // @[TBE.scala 112:26]
  wire  _GEN_1617 = _GEN_4172 | _GEN_1536; // @[TBE.scala 112:26]
  wire  _GEN_1618 = _GEN_4173 | _GEN_1537; // @[TBE.scala 112:26]
  wire  _GEN_1619 = _GEN_4174 | _GEN_1538; // @[TBE.scala 112:26]
  wire  _GEN_1620 = _GEN_4175 | _GEN_1539; // @[TBE.scala 112:26]
  wire  _GEN_1621 = _GEN_4176 | _GEN_1540; // @[TBE.scala 112:26]
  wire  _T_283 = io_write_3_bits_command == 2'h2; // @[TBE.scala 137:46]
  wire  isDealloc_3 = _T_283 & io_write_3_valid; // @[TBE.scala 137:58]
  wire  _T_155 = isDealloc_3 & finder_3_io_value_valid; // @[TBE.scala 114:31]
  wire [4:0] idxUpdate_3 = {{1'd0}, finder_3_io_value_bits}; // @[TBE.scala 73:23 TBE.scala 104:18]
  wire  _GEN_1622 = 4'h0 == idxUpdate_3[3:0] ? 1'h0 : _GEN_1525; // @[TBE.scala 115:30]
  wire  _GEN_1623 = 4'h1 == idxUpdate_3[3:0] ? 1'h0 : _GEN_1526; // @[TBE.scala 115:30]
  wire  _GEN_1624 = 4'h2 == idxUpdate_3[3:0] ? 1'h0 : _GEN_1527; // @[TBE.scala 115:30]
  wire  _GEN_1625 = 4'h3 == idxUpdate_3[3:0] ? 1'h0 : _GEN_1528; // @[TBE.scala 115:30]
  wire  _GEN_1626 = 4'h4 == idxUpdate_3[3:0] ? 1'h0 : _GEN_1529; // @[TBE.scala 115:30]
  wire  _GEN_1627 = 4'h5 == idxUpdate_3[3:0] ? 1'h0 : _GEN_1530; // @[TBE.scala 115:30]
  wire  _GEN_1628 = 4'h6 == idxUpdate_3[3:0] ? 1'h0 : _GEN_1531; // @[TBE.scala 115:30]
  wire  _GEN_1629 = 4'h7 == idxUpdate_3[3:0] ? 1'h0 : _GEN_1532; // @[TBE.scala 115:30]
  wire  _GEN_1630 = 4'h8 == idxUpdate_3[3:0] ? 1'h0 : _GEN_1533; // @[TBE.scala 115:30]
  wire  _GEN_1631 = 4'h9 == idxUpdate_3[3:0] ? 1'h0 : _GEN_1534; // @[TBE.scala 115:30]
  wire  _GEN_1632 = 4'ha == idxUpdate_3[3:0] ? 1'h0 : _GEN_1535; // @[TBE.scala 115:30]
  wire  _GEN_1633 = 4'hb == idxUpdate_3[3:0] ? 1'h0 : _GEN_1536; // @[TBE.scala 115:30]
  wire  _GEN_1634 = 4'hc == idxUpdate_3[3:0] ? 1'h0 : _GEN_1537; // @[TBE.scala 115:30]
  wire  _GEN_1635 = 4'hd == idxUpdate_3[3:0] ? 1'h0 : _GEN_1538; // @[TBE.scala 115:30]
  wire  _GEN_1636 = 4'he == idxUpdate_3[3:0] ? 1'h0 : _GEN_1539; // @[TBE.scala 115:30]
  wire  _GEN_1637 = 4'hf == idxUpdate_3[3:0] ? 1'h0 : _GEN_1540; // @[TBE.scala 115:30]
  wire [31:0] _GEN_1638 = 4'h0 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1461; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1639 = 4'h1 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1462; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1640 = 4'h2 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1463; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1641 = 4'h3 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1464; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1642 = 4'h4 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1465; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1643 = 4'h5 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1466; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1644 = 4'h6 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1467; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1645 = 4'h7 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1468; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1646 = 4'h8 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1469; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1647 = 4'h9 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1470; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1648 = 4'ha == idxUpdate_3[3:0] ? 32'h0 : _GEN_1471; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1649 = 4'hb == idxUpdate_3[3:0] ? 32'h0 : _GEN_1472; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1650 = 4'hc == idxUpdate_3[3:0] ? 32'h0 : _GEN_1473; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1651 = 4'hd == idxUpdate_3[3:0] ? 32'h0 : _GEN_1474; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1652 = 4'he == idxUpdate_3[3:0] ? 32'h0 : _GEN_1475; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1653 = 4'hf == idxUpdate_3[3:0] ? 32'h0 : _GEN_1476; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1654 = 4'h0 == idxUpdate_3[3:0] ? 3'h2 : _GEN_1477; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1655 = 4'h1 == idxUpdate_3[3:0] ? 3'h2 : _GEN_1478; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1656 = 4'h2 == idxUpdate_3[3:0] ? 3'h2 : _GEN_1479; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1657 = 4'h3 == idxUpdate_3[3:0] ? 3'h2 : _GEN_1480; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1658 = 4'h4 == idxUpdate_3[3:0] ? 3'h2 : _GEN_1481; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1659 = 4'h5 == idxUpdate_3[3:0] ? 3'h2 : _GEN_1482; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1660 = 4'h6 == idxUpdate_3[3:0] ? 3'h2 : _GEN_1483; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1661 = 4'h7 == idxUpdate_3[3:0] ? 3'h2 : _GEN_1484; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1662 = 4'h8 == idxUpdate_3[3:0] ? 3'h2 : _GEN_1485; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1663 = 4'h9 == idxUpdate_3[3:0] ? 3'h2 : _GEN_1486; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1664 = 4'ha == idxUpdate_3[3:0] ? 3'h2 : _GEN_1487; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1665 = 4'hb == idxUpdate_3[3:0] ? 3'h2 : _GEN_1488; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1666 = 4'hc == idxUpdate_3[3:0] ? 3'h2 : _GEN_1489; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1667 = 4'hd == idxUpdate_3[3:0] ? 3'h2 : _GEN_1490; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1668 = 4'he == idxUpdate_3[3:0] ? 3'h2 : _GEN_1491; // @[TBE.scala 116:31]
  wire [2:0] _GEN_1669 = 4'hf == idxUpdate_3[3:0] ? 3'h2 : _GEN_1492; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1670 = 4'h0 == idxUpdate_3[3:0] ? 2'h0 : _GEN_1493; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1671 = 4'h1 == idxUpdate_3[3:0] ? 2'h0 : _GEN_1494; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1672 = 4'h2 == idxUpdate_3[3:0] ? 2'h0 : _GEN_1495; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1673 = 4'h3 == idxUpdate_3[3:0] ? 2'h0 : _GEN_1496; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1674 = 4'h4 == idxUpdate_3[3:0] ? 2'h0 : _GEN_1497; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1675 = 4'h5 == idxUpdate_3[3:0] ? 2'h0 : _GEN_1498; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1676 = 4'h6 == idxUpdate_3[3:0] ? 2'h0 : _GEN_1499; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1677 = 4'h7 == idxUpdate_3[3:0] ? 2'h0 : _GEN_1500; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1678 = 4'h8 == idxUpdate_3[3:0] ? 2'h0 : _GEN_1501; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1679 = 4'h9 == idxUpdate_3[3:0] ? 2'h0 : _GEN_1502; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1680 = 4'ha == idxUpdate_3[3:0] ? 2'h0 : _GEN_1503; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1681 = 4'hb == idxUpdate_3[3:0] ? 2'h0 : _GEN_1504; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1682 = 4'hc == idxUpdate_3[3:0] ? 2'h0 : _GEN_1505; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1683 = 4'hd == idxUpdate_3[3:0] ? 2'h0 : _GEN_1506; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1684 = 4'he == idxUpdate_3[3:0] ? 2'h0 : _GEN_1507; // @[TBE.scala 116:31]
  wire [1:0] _GEN_1685 = 4'hf == idxUpdate_3[3:0] ? 2'h0 : _GEN_1508; // @[TBE.scala 116:31]
  wire [31:0] _GEN_1686 = 4'h0 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1509; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1687 = 4'h1 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1510; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1688 = 4'h2 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1511; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1689 = 4'h3 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1512; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1690 = 4'h4 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1513; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1691 = 4'h5 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1514; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1692 = 4'h6 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1515; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1693 = 4'h7 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1516; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1694 = 4'h8 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1517; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1695 = 4'h9 == idxUpdate_3[3:0] ? 32'h0 : _GEN_1518; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1696 = 4'ha == idxUpdate_3[3:0] ? 32'h0 : _GEN_1519; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1697 = 4'hb == idxUpdate_3[3:0] ? 32'h0 : _GEN_1520; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1698 = 4'hc == idxUpdate_3[3:0] ? 32'h0 : _GEN_1521; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1699 = 4'hd == idxUpdate_3[3:0] ? 32'h0 : _GEN_1522; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1700 = 4'he == idxUpdate_3[3:0] ? 32'h0 : _GEN_1523; // @[TBE.scala 117:29]
  wire [31:0] _GEN_1701 = 4'hf == idxUpdate_3[3:0] ? 32'h0 : _GEN_1524; // @[TBE.scala 117:29]
  wire  _T_285 = io_write_3_bits_command == 2'h3; // @[TBE.scala 138:44]
  wire  isWrite_3 = _T_285 & io_write_3_valid; // @[TBE.scala 138:55]
  wire  _T_163 = isWrite_3 & finder_3_io_value_valid; // @[TBE.scala 119:29]
  wire  _T_164 = ~io_write_3_bits_mask; // @[TBE.scala 120:35]
  wire [31:0] _GEN_1702 = 4'h0 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1461; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1703 = 4'h1 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1462; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1704 = 4'h2 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1463; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1705 = 4'h3 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1464; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1706 = 4'h4 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1465; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1707 = 4'h5 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1466; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1708 = 4'h6 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1467; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1709 = 4'h7 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1468; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1710 = 4'h8 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1469; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1711 = 4'h9 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1470; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1712 = 4'ha == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1471; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1713 = 4'hb == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1472; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1714 = 4'hc == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1473; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1715 = 4'hd == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1474; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1716 = 4'he == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1475; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1717 = 4'hf == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_fields_0 : _GEN_1476; // @[TBE.scala 121:63]
  wire [31:0] _GEN_1723 = 4'h1 == idxUpdate_3[3:0] ? TBEMemory_1_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1726 = 4'h2 == idxUpdate_3[3:0] ? TBEMemory_2_fields_0 : _GEN_1723; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1729 = 4'h3 == idxUpdate_3[3:0] ? TBEMemory_3_fields_0 : _GEN_1726; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1732 = 4'h4 == idxUpdate_3[3:0] ? TBEMemory_4_fields_0 : _GEN_1729; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1735 = 4'h5 == idxUpdate_3[3:0] ? TBEMemory_5_fields_0 : _GEN_1732; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1738 = 4'h6 == idxUpdate_3[3:0] ? TBEMemory_6_fields_0 : _GEN_1735; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1741 = 4'h7 == idxUpdate_3[3:0] ? TBEMemory_7_fields_0 : _GEN_1738; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1744 = 4'h8 == idxUpdate_3[3:0] ? TBEMemory_8_fields_0 : _GEN_1741; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1747 = 4'h9 == idxUpdate_3[3:0] ? TBEMemory_9_fields_0 : _GEN_1744; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1750 = 4'ha == idxUpdate_3[3:0] ? TBEMemory_10_fields_0 : _GEN_1747; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1753 = 4'hb == idxUpdate_3[3:0] ? TBEMemory_11_fields_0 : _GEN_1750; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1756 = 4'hc == idxUpdate_3[3:0] ? TBEMemory_12_fields_0 : _GEN_1753; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1759 = 4'hd == idxUpdate_3[3:0] ? TBEMemory_13_fields_0 : _GEN_1756; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1762 = 4'he == idxUpdate_3[3:0] ? TBEMemory_14_fields_0 : _GEN_1759; // @[TBE.scala 122:15]
  wire [31:0] _GEN_1765 = 4'hf == idxUpdate_3[3:0] ? TBEMemory_15_fields_0 : _GEN_1762; // @[TBE.scala 122:15]
  wire [2:0] _GEN_1766 = 4'h0 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1477; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1767 = 4'h1 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1478; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1768 = 4'h2 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1479; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1769 = 4'h3 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1480; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1770 = 4'h4 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1481; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1771 = 4'h5 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1482; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1772 = 4'h6 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1483; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1773 = 4'h7 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1484; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1774 = 4'h8 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1485; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1775 = 4'h9 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1486; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1776 = 4'ha == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1487; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1777 = 4'hb == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1488; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1778 = 4'hc == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1489; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1779 = 4'hd == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1490; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1780 = 4'he == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1491; // @[TBE.scala 124:37]
  wire [2:0] _GEN_1781 = 4'hf == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_way : _GEN_1492; // @[TBE.scala 124:37]
  wire [1:0] _GEN_1782 = 4'h0 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1493; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1783 = 4'h1 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1494; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1784 = 4'h2 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1495; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1785 = 4'h3 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1496; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1786 = 4'h4 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1497; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1787 = 4'h5 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1498; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1788 = 4'h6 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1499; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1789 = 4'h7 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1500; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1790 = 4'h8 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1501; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1791 = 4'h9 == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1502; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1792 = 4'ha == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1503; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1793 = 4'hb == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1504; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1794 = 4'hc == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1505; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1795 = 4'hd == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1506; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1796 = 4'he == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1507; // @[TBE.scala 125:39]
  wire [1:0] _GEN_1797 = 4'hf == idxUpdate_3[3:0] ? io_write_3_bits_inputTBE_state_state : _GEN_1508; // @[TBE.scala 125:39]
  wire [31:0] _GEN_1798 = _T_164 ? _GEN_1702 : _GEN_1461; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1799 = _T_164 ? _GEN_1703 : _GEN_1462; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1800 = _T_164 ? _GEN_1704 : _GEN_1463; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1801 = _T_164 ? _GEN_1705 : _GEN_1464; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1802 = _T_164 ? _GEN_1706 : _GEN_1465; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1803 = _T_164 ? _GEN_1707 : _GEN_1466; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1804 = _T_164 ? _GEN_1708 : _GEN_1467; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1805 = _T_164 ? _GEN_1709 : _GEN_1468; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1806 = _T_164 ? _GEN_1710 : _GEN_1469; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1807 = _T_164 ? _GEN_1711 : _GEN_1470; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1808 = _T_164 ? _GEN_1712 : _GEN_1471; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1809 = _T_164 ? _GEN_1713 : _GEN_1472; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1810 = _T_164 ? _GEN_1714 : _GEN_1473; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1811 = _T_164 ? _GEN_1715 : _GEN_1474; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1812 = _T_164 ? _GEN_1716 : _GEN_1475; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1813 = _T_164 ? _GEN_1717 : _GEN_1476; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1814 = _T_164 ? _GEN_1477 : _GEN_1766; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1815 = _T_164 ? _GEN_1478 : _GEN_1767; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1816 = _T_164 ? _GEN_1479 : _GEN_1768; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1817 = _T_164 ? _GEN_1480 : _GEN_1769; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1818 = _T_164 ? _GEN_1481 : _GEN_1770; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1819 = _T_164 ? _GEN_1482 : _GEN_1771; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1820 = _T_164 ? _GEN_1483 : _GEN_1772; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1821 = _T_164 ? _GEN_1484 : _GEN_1773; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1822 = _T_164 ? _GEN_1485 : _GEN_1774; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1823 = _T_164 ? _GEN_1486 : _GEN_1775; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1824 = _T_164 ? _GEN_1487 : _GEN_1776; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1825 = _T_164 ? _GEN_1488 : _GEN_1777; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1826 = _T_164 ? _GEN_1489 : _GEN_1778; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1827 = _T_164 ? _GEN_1490 : _GEN_1779; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1828 = _T_164 ? _GEN_1491 : _GEN_1780; // @[TBE.scala 120:53]
  wire [2:0] _GEN_1829 = _T_164 ? _GEN_1492 : _GEN_1781; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1830 = _T_164 ? _GEN_1493 : _GEN_1782; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1831 = _T_164 ? _GEN_1494 : _GEN_1783; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1832 = _T_164 ? _GEN_1495 : _GEN_1784; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1833 = _T_164 ? _GEN_1496 : _GEN_1785; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1834 = _T_164 ? _GEN_1497 : _GEN_1786; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1835 = _T_164 ? _GEN_1498 : _GEN_1787; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1836 = _T_164 ? _GEN_1499 : _GEN_1788; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1837 = _T_164 ? _GEN_1500 : _GEN_1789; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1838 = _T_164 ? _GEN_1501 : _GEN_1790; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1839 = _T_164 ? _GEN_1502 : _GEN_1791; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1840 = _T_164 ? _GEN_1503 : _GEN_1792; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1841 = _T_164 ? _GEN_1504 : _GEN_1793; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1842 = _T_164 ? _GEN_1505 : _GEN_1794; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1843 = _T_164 ? _GEN_1506 : _GEN_1795; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1844 = _T_164 ? _GEN_1507 : _GEN_1796; // @[TBE.scala 120:53]
  wire [1:0] _GEN_1845 = _T_164 ? _GEN_1508 : _GEN_1797; // @[TBE.scala 120:53]
  wire [31:0] _GEN_1846 = _T_163 ? _GEN_1798 : _GEN_1461; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1847 = _T_163 ? _GEN_1799 : _GEN_1462; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1848 = _T_163 ? _GEN_1800 : _GEN_1463; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1849 = _T_163 ? _GEN_1801 : _GEN_1464; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1850 = _T_163 ? _GEN_1802 : _GEN_1465; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1851 = _T_163 ? _GEN_1803 : _GEN_1466; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1852 = _T_163 ? _GEN_1804 : _GEN_1467; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1853 = _T_163 ? _GEN_1805 : _GEN_1468; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1854 = _T_163 ? _GEN_1806 : _GEN_1469; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1855 = _T_163 ? _GEN_1807 : _GEN_1470; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1856 = _T_163 ? _GEN_1808 : _GEN_1471; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1857 = _T_163 ? _GEN_1809 : _GEN_1472; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1858 = _T_163 ? _GEN_1810 : _GEN_1473; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1859 = _T_163 ? _GEN_1811 : _GEN_1474; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1860 = _T_163 ? _GEN_1812 : _GEN_1475; // @[TBE.scala 119:57]
  wire [31:0] _GEN_1861 = _T_163 ? _GEN_1813 : _GEN_1476; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1862 = _T_163 ? _GEN_1814 : _GEN_1477; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1863 = _T_163 ? _GEN_1815 : _GEN_1478; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1864 = _T_163 ? _GEN_1816 : _GEN_1479; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1865 = _T_163 ? _GEN_1817 : _GEN_1480; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1866 = _T_163 ? _GEN_1818 : _GEN_1481; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1867 = _T_163 ? _GEN_1819 : _GEN_1482; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1868 = _T_163 ? _GEN_1820 : _GEN_1483; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1869 = _T_163 ? _GEN_1821 : _GEN_1484; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1870 = _T_163 ? _GEN_1822 : _GEN_1485; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1871 = _T_163 ? _GEN_1823 : _GEN_1486; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1872 = _T_163 ? _GEN_1824 : _GEN_1487; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1873 = _T_163 ? _GEN_1825 : _GEN_1488; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1874 = _T_163 ? _GEN_1826 : _GEN_1489; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1875 = _T_163 ? _GEN_1827 : _GEN_1490; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1876 = _T_163 ? _GEN_1828 : _GEN_1491; // @[TBE.scala 119:57]
  wire [2:0] _GEN_1877 = _T_163 ? _GEN_1829 : _GEN_1492; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1878 = _T_163 ? _GEN_1830 : _GEN_1493; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1879 = _T_163 ? _GEN_1831 : _GEN_1494; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1880 = _T_163 ? _GEN_1832 : _GEN_1495; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1881 = _T_163 ? _GEN_1833 : _GEN_1496; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1882 = _T_163 ? _GEN_1834 : _GEN_1497; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1883 = _T_163 ? _GEN_1835 : _GEN_1498; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1884 = _T_163 ? _GEN_1836 : _GEN_1499; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1885 = _T_163 ? _GEN_1837 : _GEN_1500; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1886 = _T_163 ? _GEN_1838 : _GEN_1501; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1887 = _T_163 ? _GEN_1839 : _GEN_1502; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1888 = _T_163 ? _GEN_1840 : _GEN_1503; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1889 = _T_163 ? _GEN_1841 : _GEN_1504; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1890 = _T_163 ? _GEN_1842 : _GEN_1505; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1891 = _T_163 ? _GEN_1843 : _GEN_1506; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1892 = _T_163 ? _GEN_1844 : _GEN_1507; // @[TBE.scala 119:57]
  wire [1:0] _GEN_1893 = _T_163 ? _GEN_1845 : _GEN_1508; // @[TBE.scala 119:57]
  wire  _GEN_1894 = _T_155 ? _GEN_1622 : _GEN_1525; // @[TBE.scala 114:59]
  wire  _GEN_1895 = _T_155 ? _GEN_1623 : _GEN_1526; // @[TBE.scala 114:59]
  wire  _GEN_1896 = _T_155 ? _GEN_1624 : _GEN_1527; // @[TBE.scala 114:59]
  wire  _GEN_1897 = _T_155 ? _GEN_1625 : _GEN_1528; // @[TBE.scala 114:59]
  wire  _GEN_1898 = _T_155 ? _GEN_1626 : _GEN_1529; // @[TBE.scala 114:59]
  wire  _GEN_1899 = _T_155 ? _GEN_1627 : _GEN_1530; // @[TBE.scala 114:59]
  wire  _GEN_1900 = _T_155 ? _GEN_1628 : _GEN_1531; // @[TBE.scala 114:59]
  wire  _GEN_1901 = _T_155 ? _GEN_1629 : _GEN_1532; // @[TBE.scala 114:59]
  wire  _GEN_1902 = _T_155 ? _GEN_1630 : _GEN_1533; // @[TBE.scala 114:59]
  wire  _GEN_1903 = _T_155 ? _GEN_1631 : _GEN_1534; // @[TBE.scala 114:59]
  wire  _GEN_1904 = _T_155 ? _GEN_1632 : _GEN_1535; // @[TBE.scala 114:59]
  wire  _GEN_1905 = _T_155 ? _GEN_1633 : _GEN_1536; // @[TBE.scala 114:59]
  wire  _GEN_1906 = _T_155 ? _GEN_1634 : _GEN_1537; // @[TBE.scala 114:59]
  wire  _GEN_1907 = _T_155 ? _GEN_1635 : _GEN_1538; // @[TBE.scala 114:59]
  wire  _GEN_1908 = _T_155 ? _GEN_1636 : _GEN_1539; // @[TBE.scala 114:59]
  wire  _GEN_1909 = _T_155 ? _GEN_1637 : _GEN_1540; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1910 = _T_155 ? _GEN_1638 : _GEN_1846; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1911 = _T_155 ? _GEN_1639 : _GEN_1847; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1912 = _T_155 ? _GEN_1640 : _GEN_1848; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1913 = _T_155 ? _GEN_1641 : _GEN_1849; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1914 = _T_155 ? _GEN_1642 : _GEN_1850; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1915 = _T_155 ? _GEN_1643 : _GEN_1851; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1916 = _T_155 ? _GEN_1644 : _GEN_1852; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1917 = _T_155 ? _GEN_1645 : _GEN_1853; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1918 = _T_155 ? _GEN_1646 : _GEN_1854; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1919 = _T_155 ? _GEN_1647 : _GEN_1855; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1920 = _T_155 ? _GEN_1648 : _GEN_1856; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1921 = _T_155 ? _GEN_1649 : _GEN_1857; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1922 = _T_155 ? _GEN_1650 : _GEN_1858; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1923 = _T_155 ? _GEN_1651 : _GEN_1859; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1924 = _T_155 ? _GEN_1652 : _GEN_1860; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1925 = _T_155 ? _GEN_1653 : _GEN_1861; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1926 = _T_155 ? _GEN_1654 : _GEN_1862; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1927 = _T_155 ? _GEN_1655 : _GEN_1863; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1928 = _T_155 ? _GEN_1656 : _GEN_1864; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1929 = _T_155 ? _GEN_1657 : _GEN_1865; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1930 = _T_155 ? _GEN_1658 : _GEN_1866; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1931 = _T_155 ? _GEN_1659 : _GEN_1867; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1932 = _T_155 ? _GEN_1660 : _GEN_1868; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1933 = _T_155 ? _GEN_1661 : _GEN_1869; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1934 = _T_155 ? _GEN_1662 : _GEN_1870; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1935 = _T_155 ? _GEN_1663 : _GEN_1871; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1936 = _T_155 ? _GEN_1664 : _GEN_1872; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1937 = _T_155 ? _GEN_1665 : _GEN_1873; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1938 = _T_155 ? _GEN_1666 : _GEN_1874; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1939 = _T_155 ? _GEN_1667 : _GEN_1875; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1940 = _T_155 ? _GEN_1668 : _GEN_1876; // @[TBE.scala 114:59]
  wire [2:0] _GEN_1941 = _T_155 ? _GEN_1669 : _GEN_1877; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1942 = _T_155 ? _GEN_1670 : _GEN_1878; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1943 = _T_155 ? _GEN_1671 : _GEN_1879; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1944 = _T_155 ? _GEN_1672 : _GEN_1880; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1945 = _T_155 ? _GEN_1673 : _GEN_1881; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1946 = _T_155 ? _GEN_1674 : _GEN_1882; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1947 = _T_155 ? _GEN_1675 : _GEN_1883; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1948 = _T_155 ? _GEN_1676 : _GEN_1884; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1949 = _T_155 ? _GEN_1677 : _GEN_1885; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1950 = _T_155 ? _GEN_1678 : _GEN_1886; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1951 = _T_155 ? _GEN_1679 : _GEN_1887; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1952 = _T_155 ? _GEN_1680 : _GEN_1888; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1953 = _T_155 ? _GEN_1681 : _GEN_1889; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1954 = _T_155 ? _GEN_1682 : _GEN_1890; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1955 = _T_155 ? _GEN_1683 : _GEN_1891; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1956 = _T_155 ? _GEN_1684 : _GEN_1892; // @[TBE.scala 114:59]
  wire [1:0] _GEN_1957 = _T_155 ? _GEN_1685 : _GEN_1893; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1958 = _T_155 ? _GEN_1686 : _GEN_1509; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1959 = _T_155 ? _GEN_1687 : _GEN_1510; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1960 = _T_155 ? _GEN_1688 : _GEN_1511; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1961 = _T_155 ? _GEN_1689 : _GEN_1512; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1962 = _T_155 ? _GEN_1690 : _GEN_1513; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1963 = _T_155 ? _GEN_1691 : _GEN_1514; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1964 = _T_155 ? _GEN_1692 : _GEN_1515; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1965 = _T_155 ? _GEN_1693 : _GEN_1516; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1966 = _T_155 ? _GEN_1694 : _GEN_1517; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1967 = _T_155 ? _GEN_1695 : _GEN_1518; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1968 = _T_155 ? _GEN_1696 : _GEN_1519; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1969 = _T_155 ? _GEN_1697 : _GEN_1520; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1970 = _T_155 ? _GEN_1698 : _GEN_1521; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1971 = _T_155 ? _GEN_1699 : _GEN_1522; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1972 = _T_155 ? _GEN_1700 : _GEN_1523; // @[TBE.scala 114:59]
  wire [31:0] _GEN_1973 = _T_155 ? _GEN_1701 : _GEN_1524; // @[TBE.scala 114:59]
  wire  _T_281 = io_write_3_bits_command == 2'h1; // @[TBE.scala 136:44]
  wire  isAlloc_3 = _T_281 & io_write_3_valid; // @[TBE.scala 136:54]
  wire [31:0] _GEN_1975 = isAlloc_3 ? _GEN_1542 : _GEN_1910; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1976 = isAlloc_3 ? _GEN_1543 : _GEN_1911; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1977 = isAlloc_3 ? _GEN_1544 : _GEN_1912; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1978 = isAlloc_3 ? _GEN_1545 : _GEN_1913; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1979 = isAlloc_3 ? _GEN_1546 : _GEN_1914; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1980 = isAlloc_3 ? _GEN_1547 : _GEN_1915; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1981 = isAlloc_3 ? _GEN_1548 : _GEN_1916; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1982 = isAlloc_3 ? _GEN_1549 : _GEN_1917; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1983 = isAlloc_3 ? _GEN_1550 : _GEN_1918; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1984 = isAlloc_3 ? _GEN_1551 : _GEN_1919; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1985 = isAlloc_3 ? _GEN_1552 : _GEN_1920; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1986 = isAlloc_3 ? _GEN_1553 : _GEN_1921; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1987 = isAlloc_3 ? _GEN_1554 : _GEN_1922; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1988 = isAlloc_3 ? _GEN_1555 : _GEN_1923; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1989 = isAlloc_3 ? _GEN_1556 : _GEN_1924; // @[TBE.scala 109:24]
  wire [31:0] _GEN_1990 = isAlloc_3 ? _GEN_1557 : _GEN_1925; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1991 = isAlloc_3 ? _GEN_1558 : _GEN_1926; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1992 = isAlloc_3 ? _GEN_1559 : _GEN_1927; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1993 = isAlloc_3 ? _GEN_1560 : _GEN_1928; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1994 = isAlloc_3 ? _GEN_1561 : _GEN_1929; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1995 = isAlloc_3 ? _GEN_1562 : _GEN_1930; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1996 = isAlloc_3 ? _GEN_1563 : _GEN_1931; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1997 = isAlloc_3 ? _GEN_1564 : _GEN_1932; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1998 = isAlloc_3 ? _GEN_1565 : _GEN_1933; // @[TBE.scala 109:24]
  wire [2:0] _GEN_1999 = isAlloc_3 ? _GEN_1566 : _GEN_1934; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2000 = isAlloc_3 ? _GEN_1567 : _GEN_1935; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2001 = isAlloc_3 ? _GEN_1568 : _GEN_1936; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2002 = isAlloc_3 ? _GEN_1569 : _GEN_1937; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2003 = isAlloc_3 ? _GEN_1570 : _GEN_1938; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2004 = isAlloc_3 ? _GEN_1571 : _GEN_1939; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2005 = isAlloc_3 ? _GEN_1572 : _GEN_1940; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2006 = isAlloc_3 ? _GEN_1573 : _GEN_1941; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2007 = isAlloc_3 ? _GEN_1574 : _GEN_1942; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2008 = isAlloc_3 ? _GEN_1575 : _GEN_1943; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2009 = isAlloc_3 ? _GEN_1576 : _GEN_1944; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2010 = isAlloc_3 ? _GEN_1577 : _GEN_1945; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2011 = isAlloc_3 ? _GEN_1578 : _GEN_1946; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2012 = isAlloc_3 ? _GEN_1579 : _GEN_1947; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2013 = isAlloc_3 ? _GEN_1580 : _GEN_1948; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2014 = isAlloc_3 ? _GEN_1581 : _GEN_1949; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2015 = isAlloc_3 ? _GEN_1582 : _GEN_1950; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2016 = isAlloc_3 ? _GEN_1583 : _GEN_1951; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2017 = isAlloc_3 ? _GEN_1584 : _GEN_1952; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2018 = isAlloc_3 ? _GEN_1585 : _GEN_1953; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2019 = isAlloc_3 ? _GEN_1586 : _GEN_1954; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2020 = isAlloc_3 ? _GEN_1587 : _GEN_1955; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2021 = isAlloc_3 ? _GEN_1588 : _GEN_1956; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2022 = isAlloc_3 ? _GEN_1589 : _GEN_1957; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2023 = isAlloc_3 ? _GEN_1590 : _GEN_1958; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2024 = isAlloc_3 ? _GEN_1591 : _GEN_1959; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2025 = isAlloc_3 ? _GEN_1592 : _GEN_1960; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2026 = isAlloc_3 ? _GEN_1593 : _GEN_1961; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2027 = isAlloc_3 ? _GEN_1594 : _GEN_1962; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2028 = isAlloc_3 ? _GEN_1595 : _GEN_1963; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2029 = isAlloc_3 ? _GEN_1596 : _GEN_1964; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2030 = isAlloc_3 ? _GEN_1597 : _GEN_1965; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2031 = isAlloc_3 ? _GEN_1598 : _GEN_1966; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2032 = isAlloc_3 ? _GEN_1599 : _GEN_1967; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2033 = isAlloc_3 ? _GEN_1600 : _GEN_1968; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2034 = isAlloc_3 ? _GEN_1601 : _GEN_1969; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2035 = isAlloc_3 ? _GEN_1602 : _GEN_1970; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2036 = isAlloc_3 ? _GEN_1603 : _GEN_1971; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2037 = isAlloc_3 ? _GEN_1604 : _GEN_1972; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2038 = isAlloc_3 ? _GEN_1605 : _GEN_1973; // @[TBE.scala 109:24]
  wire  _GEN_2039 = isAlloc_3 ? _GEN_1606 : _GEN_1894; // @[TBE.scala 109:24]
  wire  _GEN_2040 = isAlloc_3 ? _GEN_1607 : _GEN_1895; // @[TBE.scala 109:24]
  wire  _GEN_2041 = isAlloc_3 ? _GEN_1608 : _GEN_1896; // @[TBE.scala 109:24]
  wire  _GEN_2042 = isAlloc_3 ? _GEN_1609 : _GEN_1897; // @[TBE.scala 109:24]
  wire  _GEN_2043 = isAlloc_3 ? _GEN_1610 : _GEN_1898; // @[TBE.scala 109:24]
  wire  _GEN_2044 = isAlloc_3 ? _GEN_1611 : _GEN_1899; // @[TBE.scala 109:24]
  wire  _GEN_2045 = isAlloc_3 ? _GEN_1612 : _GEN_1900; // @[TBE.scala 109:24]
  wire  _GEN_2046 = isAlloc_3 ? _GEN_1613 : _GEN_1901; // @[TBE.scala 109:24]
  wire  _GEN_2047 = isAlloc_3 ? _GEN_1614 : _GEN_1902; // @[TBE.scala 109:24]
  wire  _GEN_2048 = isAlloc_3 ? _GEN_1615 : _GEN_1903; // @[TBE.scala 109:24]
  wire  _GEN_2049 = isAlloc_3 ? _GEN_1616 : _GEN_1904; // @[TBE.scala 109:24]
  wire  _GEN_2050 = isAlloc_3 ? _GEN_1617 : _GEN_1905; // @[TBE.scala 109:24]
  wire  _GEN_2051 = isAlloc_3 ? _GEN_1618 : _GEN_1906; // @[TBE.scala 109:24]
  wire  _GEN_2052 = isAlloc_3 ? _GEN_1619 : _GEN_1907; // @[TBE.scala 109:24]
  wire  _GEN_2053 = isAlloc_3 ? _GEN_1620 : _GEN_1908; // @[TBE.scala 109:24]
  wire  _GEN_2054 = isAlloc_3 ? _GEN_1621 : _GEN_1909; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2056 = 4'h0 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1975; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2057 = 4'h1 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1976; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2058 = 4'h2 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1977; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2059 = 4'h3 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1978; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2060 = 4'h4 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1979; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2061 = 4'h5 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1980; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2062 = 4'h6 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1981; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2063 = 4'h7 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1982; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2064 = 4'h8 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1983; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2065 = 4'h9 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1984; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2066 = 4'ha == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1985; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2067 = 4'hb == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1986; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2068 = 4'hc == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1987; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2069 = 4'hd == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1988; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2070 = 4'he == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1989; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2071 = 4'hf == idxAlloc[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1990; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2072 = 4'h0 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1991; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2073 = 4'h1 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1992; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2074 = 4'h2 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1993; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2075 = 4'h3 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1994; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2076 = 4'h4 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1995; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2077 = 4'h5 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1996; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2078 = 4'h6 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1997; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2079 = 4'h7 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1998; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2080 = 4'h8 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1999; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2081 = 4'h9 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2000; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2082 = 4'ha == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2001; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2083 = 4'hb == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2002; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2084 = 4'hc == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2003; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2085 = 4'hd == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2004; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2086 = 4'he == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2005; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2087 = 4'hf == idxAlloc[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2006; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2088 = 4'h0 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2007; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2089 = 4'h1 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2008; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2090 = 4'h2 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2009; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2091 = 4'h3 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2010; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2092 = 4'h4 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2011; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2093 = 4'h5 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2012; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2094 = 4'h6 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2013; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2095 = 4'h7 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2014; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2096 = 4'h8 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2015; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2097 = 4'h9 == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2016; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2098 = 4'ha == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2017; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2099 = 4'hb == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2018; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2100 = 4'hc == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2019; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2101 = 4'hd == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2020; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2102 = 4'he == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2021; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2103 = 4'hf == idxAlloc[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2022; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2104 = 4'h0 == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2023; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2105 = 4'h1 == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2024; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2106 = 4'h2 == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2025; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2107 = 4'h3 == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2026; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2108 = 4'h4 == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2027; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2109 = 4'h5 == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2028; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2110 = 4'h6 == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2029; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2111 = 4'h7 == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2030; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2112 = 4'h8 == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2031; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2113 = 4'h9 == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2032; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2114 = 4'ha == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2033; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2115 = 4'hb == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2034; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2116 = 4'hc == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2035; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2117 = 4'hd == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2036; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2118 = 4'he == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2037; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2119 = 4'hf == idxAlloc[3:0] ? io_write_4_bits_addr[31:0] : _GEN_2038; // @[TBE.scala 111:25]
  wire  _GEN_2120 = _GEN_4161 | _GEN_2039; // @[TBE.scala 112:26]
  wire  _GEN_2121 = _GEN_4162 | _GEN_2040; // @[TBE.scala 112:26]
  wire  _GEN_2122 = _GEN_4163 | _GEN_2041; // @[TBE.scala 112:26]
  wire  _GEN_2123 = _GEN_4164 | _GEN_2042; // @[TBE.scala 112:26]
  wire  _GEN_2124 = _GEN_4165 | _GEN_2043; // @[TBE.scala 112:26]
  wire  _GEN_2125 = _GEN_4166 | _GEN_2044; // @[TBE.scala 112:26]
  wire  _GEN_2126 = _GEN_4167 | _GEN_2045; // @[TBE.scala 112:26]
  wire  _GEN_2127 = _GEN_4168 | _GEN_2046; // @[TBE.scala 112:26]
  wire  _GEN_2128 = _GEN_4169 | _GEN_2047; // @[TBE.scala 112:26]
  wire  _GEN_2129 = _GEN_4170 | _GEN_2048; // @[TBE.scala 112:26]
  wire  _GEN_2130 = _GEN_4171 | _GEN_2049; // @[TBE.scala 112:26]
  wire  _GEN_2131 = _GEN_4172 | _GEN_2050; // @[TBE.scala 112:26]
  wire  _GEN_2132 = _GEN_4173 | _GEN_2051; // @[TBE.scala 112:26]
  wire  _GEN_2133 = _GEN_4174 | _GEN_2052; // @[TBE.scala 112:26]
  wire  _GEN_2134 = _GEN_4175 | _GEN_2053; // @[TBE.scala 112:26]
  wire  _GEN_2135 = _GEN_4176 | _GEN_2054; // @[TBE.scala 112:26]
  wire  _T_289 = io_write_4_bits_command == 2'h2; // @[TBE.scala 137:46]
  wire  isDealloc_4 = _T_289 & io_write_4_valid; // @[TBE.scala 137:58]
  wire  _T_177 = isDealloc_4 & finder_4_io_value_valid; // @[TBE.scala 114:31]
  wire [4:0] idxUpdate_4 = {{1'd0}, finder_4_io_value_bits}; // @[TBE.scala 73:23 TBE.scala 104:18]
  wire  _GEN_2136 = 4'h0 == idxUpdate_4[3:0] ? 1'h0 : _GEN_2039; // @[TBE.scala 115:30]
  wire  _GEN_2137 = 4'h1 == idxUpdate_4[3:0] ? 1'h0 : _GEN_2040; // @[TBE.scala 115:30]
  wire  _GEN_2138 = 4'h2 == idxUpdate_4[3:0] ? 1'h0 : _GEN_2041; // @[TBE.scala 115:30]
  wire  _GEN_2139 = 4'h3 == idxUpdate_4[3:0] ? 1'h0 : _GEN_2042; // @[TBE.scala 115:30]
  wire  _GEN_2140 = 4'h4 == idxUpdate_4[3:0] ? 1'h0 : _GEN_2043; // @[TBE.scala 115:30]
  wire  _GEN_2141 = 4'h5 == idxUpdate_4[3:0] ? 1'h0 : _GEN_2044; // @[TBE.scala 115:30]
  wire  _GEN_2142 = 4'h6 == idxUpdate_4[3:0] ? 1'h0 : _GEN_2045; // @[TBE.scala 115:30]
  wire  _GEN_2143 = 4'h7 == idxUpdate_4[3:0] ? 1'h0 : _GEN_2046; // @[TBE.scala 115:30]
  wire  _GEN_2144 = 4'h8 == idxUpdate_4[3:0] ? 1'h0 : _GEN_2047; // @[TBE.scala 115:30]
  wire  _GEN_2145 = 4'h9 == idxUpdate_4[3:0] ? 1'h0 : _GEN_2048; // @[TBE.scala 115:30]
  wire  _GEN_2146 = 4'ha == idxUpdate_4[3:0] ? 1'h0 : _GEN_2049; // @[TBE.scala 115:30]
  wire  _GEN_2147 = 4'hb == idxUpdate_4[3:0] ? 1'h0 : _GEN_2050; // @[TBE.scala 115:30]
  wire  _GEN_2148 = 4'hc == idxUpdate_4[3:0] ? 1'h0 : _GEN_2051; // @[TBE.scala 115:30]
  wire  _GEN_2149 = 4'hd == idxUpdate_4[3:0] ? 1'h0 : _GEN_2052; // @[TBE.scala 115:30]
  wire  _GEN_2150 = 4'he == idxUpdate_4[3:0] ? 1'h0 : _GEN_2053; // @[TBE.scala 115:30]
  wire  _GEN_2151 = 4'hf == idxUpdate_4[3:0] ? 1'h0 : _GEN_2054; // @[TBE.scala 115:30]
  wire [31:0] _GEN_2152 = 4'h0 == idxUpdate_4[3:0] ? 32'h0 : _GEN_1975; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2153 = 4'h1 == idxUpdate_4[3:0] ? 32'h0 : _GEN_1976; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2154 = 4'h2 == idxUpdate_4[3:0] ? 32'h0 : _GEN_1977; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2155 = 4'h3 == idxUpdate_4[3:0] ? 32'h0 : _GEN_1978; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2156 = 4'h4 == idxUpdate_4[3:0] ? 32'h0 : _GEN_1979; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2157 = 4'h5 == idxUpdate_4[3:0] ? 32'h0 : _GEN_1980; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2158 = 4'h6 == idxUpdate_4[3:0] ? 32'h0 : _GEN_1981; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2159 = 4'h7 == idxUpdate_4[3:0] ? 32'h0 : _GEN_1982; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2160 = 4'h8 == idxUpdate_4[3:0] ? 32'h0 : _GEN_1983; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2161 = 4'h9 == idxUpdate_4[3:0] ? 32'h0 : _GEN_1984; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2162 = 4'ha == idxUpdate_4[3:0] ? 32'h0 : _GEN_1985; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2163 = 4'hb == idxUpdate_4[3:0] ? 32'h0 : _GEN_1986; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2164 = 4'hc == idxUpdate_4[3:0] ? 32'h0 : _GEN_1987; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2165 = 4'hd == idxUpdate_4[3:0] ? 32'h0 : _GEN_1988; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2166 = 4'he == idxUpdate_4[3:0] ? 32'h0 : _GEN_1989; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2167 = 4'hf == idxUpdate_4[3:0] ? 32'h0 : _GEN_1990; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2168 = 4'h0 == idxUpdate_4[3:0] ? 3'h2 : _GEN_1991; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2169 = 4'h1 == idxUpdate_4[3:0] ? 3'h2 : _GEN_1992; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2170 = 4'h2 == idxUpdate_4[3:0] ? 3'h2 : _GEN_1993; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2171 = 4'h3 == idxUpdate_4[3:0] ? 3'h2 : _GEN_1994; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2172 = 4'h4 == idxUpdate_4[3:0] ? 3'h2 : _GEN_1995; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2173 = 4'h5 == idxUpdate_4[3:0] ? 3'h2 : _GEN_1996; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2174 = 4'h6 == idxUpdate_4[3:0] ? 3'h2 : _GEN_1997; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2175 = 4'h7 == idxUpdate_4[3:0] ? 3'h2 : _GEN_1998; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2176 = 4'h8 == idxUpdate_4[3:0] ? 3'h2 : _GEN_1999; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2177 = 4'h9 == idxUpdate_4[3:0] ? 3'h2 : _GEN_2000; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2178 = 4'ha == idxUpdate_4[3:0] ? 3'h2 : _GEN_2001; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2179 = 4'hb == idxUpdate_4[3:0] ? 3'h2 : _GEN_2002; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2180 = 4'hc == idxUpdate_4[3:0] ? 3'h2 : _GEN_2003; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2181 = 4'hd == idxUpdate_4[3:0] ? 3'h2 : _GEN_2004; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2182 = 4'he == idxUpdate_4[3:0] ? 3'h2 : _GEN_2005; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2183 = 4'hf == idxUpdate_4[3:0] ? 3'h2 : _GEN_2006; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2184 = 4'h0 == idxUpdate_4[3:0] ? 2'h0 : _GEN_2007; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2185 = 4'h1 == idxUpdate_4[3:0] ? 2'h0 : _GEN_2008; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2186 = 4'h2 == idxUpdate_4[3:0] ? 2'h0 : _GEN_2009; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2187 = 4'h3 == idxUpdate_4[3:0] ? 2'h0 : _GEN_2010; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2188 = 4'h4 == idxUpdate_4[3:0] ? 2'h0 : _GEN_2011; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2189 = 4'h5 == idxUpdate_4[3:0] ? 2'h0 : _GEN_2012; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2190 = 4'h6 == idxUpdate_4[3:0] ? 2'h0 : _GEN_2013; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2191 = 4'h7 == idxUpdate_4[3:0] ? 2'h0 : _GEN_2014; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2192 = 4'h8 == idxUpdate_4[3:0] ? 2'h0 : _GEN_2015; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2193 = 4'h9 == idxUpdate_4[3:0] ? 2'h0 : _GEN_2016; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2194 = 4'ha == idxUpdate_4[3:0] ? 2'h0 : _GEN_2017; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2195 = 4'hb == idxUpdate_4[3:0] ? 2'h0 : _GEN_2018; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2196 = 4'hc == idxUpdate_4[3:0] ? 2'h0 : _GEN_2019; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2197 = 4'hd == idxUpdate_4[3:0] ? 2'h0 : _GEN_2020; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2198 = 4'he == idxUpdate_4[3:0] ? 2'h0 : _GEN_2021; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2199 = 4'hf == idxUpdate_4[3:0] ? 2'h0 : _GEN_2022; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2200 = 4'h0 == idxUpdate_4[3:0] ? 32'h0 : _GEN_2023; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2201 = 4'h1 == idxUpdate_4[3:0] ? 32'h0 : _GEN_2024; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2202 = 4'h2 == idxUpdate_4[3:0] ? 32'h0 : _GEN_2025; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2203 = 4'h3 == idxUpdate_4[3:0] ? 32'h0 : _GEN_2026; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2204 = 4'h4 == idxUpdate_4[3:0] ? 32'h0 : _GEN_2027; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2205 = 4'h5 == idxUpdate_4[3:0] ? 32'h0 : _GEN_2028; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2206 = 4'h6 == idxUpdate_4[3:0] ? 32'h0 : _GEN_2029; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2207 = 4'h7 == idxUpdate_4[3:0] ? 32'h0 : _GEN_2030; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2208 = 4'h8 == idxUpdate_4[3:0] ? 32'h0 : _GEN_2031; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2209 = 4'h9 == idxUpdate_4[3:0] ? 32'h0 : _GEN_2032; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2210 = 4'ha == idxUpdate_4[3:0] ? 32'h0 : _GEN_2033; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2211 = 4'hb == idxUpdate_4[3:0] ? 32'h0 : _GEN_2034; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2212 = 4'hc == idxUpdate_4[3:0] ? 32'h0 : _GEN_2035; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2213 = 4'hd == idxUpdate_4[3:0] ? 32'h0 : _GEN_2036; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2214 = 4'he == idxUpdate_4[3:0] ? 32'h0 : _GEN_2037; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2215 = 4'hf == idxUpdate_4[3:0] ? 32'h0 : _GEN_2038; // @[TBE.scala 117:29]
  wire  _T_291 = io_write_4_bits_command == 2'h3; // @[TBE.scala 138:44]
  wire  isWrite_4 = _T_291 & io_write_4_valid; // @[TBE.scala 138:55]
  wire  _T_185 = isWrite_4 & finder_4_io_value_valid; // @[TBE.scala 119:29]
  wire  _T_186 = ~io_write_4_bits_mask; // @[TBE.scala 120:35]
  wire [31:0] _GEN_2216 = 4'h0 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1975; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2217 = 4'h1 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1976; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2218 = 4'h2 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1977; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2219 = 4'h3 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1978; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2220 = 4'h4 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1979; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2221 = 4'h5 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1980; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2222 = 4'h6 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1981; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2223 = 4'h7 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1982; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2224 = 4'h8 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1983; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2225 = 4'h9 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1984; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2226 = 4'ha == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1985; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2227 = 4'hb == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1986; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2228 = 4'hc == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1987; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2229 = 4'hd == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1988; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2230 = 4'he == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1989; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2231 = 4'hf == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_fields_0 : _GEN_1990; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2237 = 4'h1 == idxUpdate_4[3:0] ? TBEMemory_1_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2240 = 4'h2 == idxUpdate_4[3:0] ? TBEMemory_2_fields_0 : _GEN_2237; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2243 = 4'h3 == idxUpdate_4[3:0] ? TBEMemory_3_fields_0 : _GEN_2240; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2246 = 4'h4 == idxUpdate_4[3:0] ? TBEMemory_4_fields_0 : _GEN_2243; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2249 = 4'h5 == idxUpdate_4[3:0] ? TBEMemory_5_fields_0 : _GEN_2246; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2252 = 4'h6 == idxUpdate_4[3:0] ? TBEMemory_6_fields_0 : _GEN_2249; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2255 = 4'h7 == idxUpdate_4[3:0] ? TBEMemory_7_fields_0 : _GEN_2252; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2258 = 4'h8 == idxUpdate_4[3:0] ? TBEMemory_8_fields_0 : _GEN_2255; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2261 = 4'h9 == idxUpdate_4[3:0] ? TBEMemory_9_fields_0 : _GEN_2258; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2264 = 4'ha == idxUpdate_4[3:0] ? TBEMemory_10_fields_0 : _GEN_2261; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2267 = 4'hb == idxUpdate_4[3:0] ? TBEMemory_11_fields_0 : _GEN_2264; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2270 = 4'hc == idxUpdate_4[3:0] ? TBEMemory_12_fields_0 : _GEN_2267; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2273 = 4'hd == idxUpdate_4[3:0] ? TBEMemory_13_fields_0 : _GEN_2270; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2276 = 4'he == idxUpdate_4[3:0] ? TBEMemory_14_fields_0 : _GEN_2273; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2279 = 4'hf == idxUpdate_4[3:0] ? TBEMemory_15_fields_0 : _GEN_2276; // @[TBE.scala 122:15]
  wire [2:0] _GEN_2280 = 4'h0 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1991; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2281 = 4'h1 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1992; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2282 = 4'h2 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1993; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2283 = 4'h3 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1994; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2284 = 4'h4 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1995; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2285 = 4'h5 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1996; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2286 = 4'h6 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1997; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2287 = 4'h7 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1998; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2288 = 4'h8 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_1999; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2289 = 4'h9 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2000; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2290 = 4'ha == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2001; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2291 = 4'hb == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2002; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2292 = 4'hc == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2003; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2293 = 4'hd == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2004; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2294 = 4'he == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2005; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2295 = 4'hf == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_way : _GEN_2006; // @[TBE.scala 124:37]
  wire [1:0] _GEN_2296 = 4'h0 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2007; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2297 = 4'h1 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2008; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2298 = 4'h2 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2009; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2299 = 4'h3 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2010; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2300 = 4'h4 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2011; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2301 = 4'h5 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2012; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2302 = 4'h6 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2013; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2303 = 4'h7 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2014; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2304 = 4'h8 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2015; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2305 = 4'h9 == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2016; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2306 = 4'ha == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2017; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2307 = 4'hb == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2018; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2308 = 4'hc == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2019; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2309 = 4'hd == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2020; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2310 = 4'he == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2021; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2311 = 4'hf == idxUpdate_4[3:0] ? io_write_4_bits_inputTBE_state_state : _GEN_2022; // @[TBE.scala 125:39]
  wire [31:0] _GEN_2312 = _T_186 ? _GEN_2216 : _GEN_1975; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2313 = _T_186 ? _GEN_2217 : _GEN_1976; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2314 = _T_186 ? _GEN_2218 : _GEN_1977; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2315 = _T_186 ? _GEN_2219 : _GEN_1978; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2316 = _T_186 ? _GEN_2220 : _GEN_1979; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2317 = _T_186 ? _GEN_2221 : _GEN_1980; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2318 = _T_186 ? _GEN_2222 : _GEN_1981; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2319 = _T_186 ? _GEN_2223 : _GEN_1982; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2320 = _T_186 ? _GEN_2224 : _GEN_1983; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2321 = _T_186 ? _GEN_2225 : _GEN_1984; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2322 = _T_186 ? _GEN_2226 : _GEN_1985; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2323 = _T_186 ? _GEN_2227 : _GEN_1986; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2324 = _T_186 ? _GEN_2228 : _GEN_1987; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2325 = _T_186 ? _GEN_2229 : _GEN_1988; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2326 = _T_186 ? _GEN_2230 : _GEN_1989; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2327 = _T_186 ? _GEN_2231 : _GEN_1990; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2328 = _T_186 ? _GEN_1991 : _GEN_2280; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2329 = _T_186 ? _GEN_1992 : _GEN_2281; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2330 = _T_186 ? _GEN_1993 : _GEN_2282; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2331 = _T_186 ? _GEN_1994 : _GEN_2283; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2332 = _T_186 ? _GEN_1995 : _GEN_2284; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2333 = _T_186 ? _GEN_1996 : _GEN_2285; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2334 = _T_186 ? _GEN_1997 : _GEN_2286; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2335 = _T_186 ? _GEN_1998 : _GEN_2287; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2336 = _T_186 ? _GEN_1999 : _GEN_2288; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2337 = _T_186 ? _GEN_2000 : _GEN_2289; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2338 = _T_186 ? _GEN_2001 : _GEN_2290; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2339 = _T_186 ? _GEN_2002 : _GEN_2291; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2340 = _T_186 ? _GEN_2003 : _GEN_2292; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2341 = _T_186 ? _GEN_2004 : _GEN_2293; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2342 = _T_186 ? _GEN_2005 : _GEN_2294; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2343 = _T_186 ? _GEN_2006 : _GEN_2295; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2344 = _T_186 ? _GEN_2007 : _GEN_2296; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2345 = _T_186 ? _GEN_2008 : _GEN_2297; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2346 = _T_186 ? _GEN_2009 : _GEN_2298; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2347 = _T_186 ? _GEN_2010 : _GEN_2299; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2348 = _T_186 ? _GEN_2011 : _GEN_2300; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2349 = _T_186 ? _GEN_2012 : _GEN_2301; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2350 = _T_186 ? _GEN_2013 : _GEN_2302; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2351 = _T_186 ? _GEN_2014 : _GEN_2303; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2352 = _T_186 ? _GEN_2015 : _GEN_2304; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2353 = _T_186 ? _GEN_2016 : _GEN_2305; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2354 = _T_186 ? _GEN_2017 : _GEN_2306; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2355 = _T_186 ? _GEN_2018 : _GEN_2307; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2356 = _T_186 ? _GEN_2019 : _GEN_2308; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2357 = _T_186 ? _GEN_2020 : _GEN_2309; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2358 = _T_186 ? _GEN_2021 : _GEN_2310; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2359 = _T_186 ? _GEN_2022 : _GEN_2311; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2360 = _T_185 ? _GEN_2312 : _GEN_1975; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2361 = _T_185 ? _GEN_2313 : _GEN_1976; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2362 = _T_185 ? _GEN_2314 : _GEN_1977; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2363 = _T_185 ? _GEN_2315 : _GEN_1978; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2364 = _T_185 ? _GEN_2316 : _GEN_1979; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2365 = _T_185 ? _GEN_2317 : _GEN_1980; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2366 = _T_185 ? _GEN_2318 : _GEN_1981; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2367 = _T_185 ? _GEN_2319 : _GEN_1982; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2368 = _T_185 ? _GEN_2320 : _GEN_1983; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2369 = _T_185 ? _GEN_2321 : _GEN_1984; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2370 = _T_185 ? _GEN_2322 : _GEN_1985; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2371 = _T_185 ? _GEN_2323 : _GEN_1986; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2372 = _T_185 ? _GEN_2324 : _GEN_1987; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2373 = _T_185 ? _GEN_2325 : _GEN_1988; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2374 = _T_185 ? _GEN_2326 : _GEN_1989; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2375 = _T_185 ? _GEN_2327 : _GEN_1990; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2376 = _T_185 ? _GEN_2328 : _GEN_1991; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2377 = _T_185 ? _GEN_2329 : _GEN_1992; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2378 = _T_185 ? _GEN_2330 : _GEN_1993; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2379 = _T_185 ? _GEN_2331 : _GEN_1994; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2380 = _T_185 ? _GEN_2332 : _GEN_1995; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2381 = _T_185 ? _GEN_2333 : _GEN_1996; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2382 = _T_185 ? _GEN_2334 : _GEN_1997; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2383 = _T_185 ? _GEN_2335 : _GEN_1998; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2384 = _T_185 ? _GEN_2336 : _GEN_1999; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2385 = _T_185 ? _GEN_2337 : _GEN_2000; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2386 = _T_185 ? _GEN_2338 : _GEN_2001; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2387 = _T_185 ? _GEN_2339 : _GEN_2002; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2388 = _T_185 ? _GEN_2340 : _GEN_2003; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2389 = _T_185 ? _GEN_2341 : _GEN_2004; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2390 = _T_185 ? _GEN_2342 : _GEN_2005; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2391 = _T_185 ? _GEN_2343 : _GEN_2006; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2392 = _T_185 ? _GEN_2344 : _GEN_2007; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2393 = _T_185 ? _GEN_2345 : _GEN_2008; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2394 = _T_185 ? _GEN_2346 : _GEN_2009; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2395 = _T_185 ? _GEN_2347 : _GEN_2010; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2396 = _T_185 ? _GEN_2348 : _GEN_2011; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2397 = _T_185 ? _GEN_2349 : _GEN_2012; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2398 = _T_185 ? _GEN_2350 : _GEN_2013; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2399 = _T_185 ? _GEN_2351 : _GEN_2014; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2400 = _T_185 ? _GEN_2352 : _GEN_2015; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2401 = _T_185 ? _GEN_2353 : _GEN_2016; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2402 = _T_185 ? _GEN_2354 : _GEN_2017; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2403 = _T_185 ? _GEN_2355 : _GEN_2018; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2404 = _T_185 ? _GEN_2356 : _GEN_2019; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2405 = _T_185 ? _GEN_2357 : _GEN_2020; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2406 = _T_185 ? _GEN_2358 : _GEN_2021; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2407 = _T_185 ? _GEN_2359 : _GEN_2022; // @[TBE.scala 119:57]
  wire  _GEN_2408 = _T_177 ? _GEN_2136 : _GEN_2039; // @[TBE.scala 114:59]
  wire  _GEN_2409 = _T_177 ? _GEN_2137 : _GEN_2040; // @[TBE.scala 114:59]
  wire  _GEN_2410 = _T_177 ? _GEN_2138 : _GEN_2041; // @[TBE.scala 114:59]
  wire  _GEN_2411 = _T_177 ? _GEN_2139 : _GEN_2042; // @[TBE.scala 114:59]
  wire  _GEN_2412 = _T_177 ? _GEN_2140 : _GEN_2043; // @[TBE.scala 114:59]
  wire  _GEN_2413 = _T_177 ? _GEN_2141 : _GEN_2044; // @[TBE.scala 114:59]
  wire  _GEN_2414 = _T_177 ? _GEN_2142 : _GEN_2045; // @[TBE.scala 114:59]
  wire  _GEN_2415 = _T_177 ? _GEN_2143 : _GEN_2046; // @[TBE.scala 114:59]
  wire  _GEN_2416 = _T_177 ? _GEN_2144 : _GEN_2047; // @[TBE.scala 114:59]
  wire  _GEN_2417 = _T_177 ? _GEN_2145 : _GEN_2048; // @[TBE.scala 114:59]
  wire  _GEN_2418 = _T_177 ? _GEN_2146 : _GEN_2049; // @[TBE.scala 114:59]
  wire  _GEN_2419 = _T_177 ? _GEN_2147 : _GEN_2050; // @[TBE.scala 114:59]
  wire  _GEN_2420 = _T_177 ? _GEN_2148 : _GEN_2051; // @[TBE.scala 114:59]
  wire  _GEN_2421 = _T_177 ? _GEN_2149 : _GEN_2052; // @[TBE.scala 114:59]
  wire  _GEN_2422 = _T_177 ? _GEN_2150 : _GEN_2053; // @[TBE.scala 114:59]
  wire  _GEN_2423 = _T_177 ? _GEN_2151 : _GEN_2054; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2424 = _T_177 ? _GEN_2152 : _GEN_2360; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2425 = _T_177 ? _GEN_2153 : _GEN_2361; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2426 = _T_177 ? _GEN_2154 : _GEN_2362; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2427 = _T_177 ? _GEN_2155 : _GEN_2363; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2428 = _T_177 ? _GEN_2156 : _GEN_2364; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2429 = _T_177 ? _GEN_2157 : _GEN_2365; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2430 = _T_177 ? _GEN_2158 : _GEN_2366; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2431 = _T_177 ? _GEN_2159 : _GEN_2367; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2432 = _T_177 ? _GEN_2160 : _GEN_2368; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2433 = _T_177 ? _GEN_2161 : _GEN_2369; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2434 = _T_177 ? _GEN_2162 : _GEN_2370; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2435 = _T_177 ? _GEN_2163 : _GEN_2371; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2436 = _T_177 ? _GEN_2164 : _GEN_2372; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2437 = _T_177 ? _GEN_2165 : _GEN_2373; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2438 = _T_177 ? _GEN_2166 : _GEN_2374; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2439 = _T_177 ? _GEN_2167 : _GEN_2375; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2440 = _T_177 ? _GEN_2168 : _GEN_2376; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2441 = _T_177 ? _GEN_2169 : _GEN_2377; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2442 = _T_177 ? _GEN_2170 : _GEN_2378; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2443 = _T_177 ? _GEN_2171 : _GEN_2379; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2444 = _T_177 ? _GEN_2172 : _GEN_2380; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2445 = _T_177 ? _GEN_2173 : _GEN_2381; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2446 = _T_177 ? _GEN_2174 : _GEN_2382; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2447 = _T_177 ? _GEN_2175 : _GEN_2383; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2448 = _T_177 ? _GEN_2176 : _GEN_2384; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2449 = _T_177 ? _GEN_2177 : _GEN_2385; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2450 = _T_177 ? _GEN_2178 : _GEN_2386; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2451 = _T_177 ? _GEN_2179 : _GEN_2387; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2452 = _T_177 ? _GEN_2180 : _GEN_2388; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2453 = _T_177 ? _GEN_2181 : _GEN_2389; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2454 = _T_177 ? _GEN_2182 : _GEN_2390; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2455 = _T_177 ? _GEN_2183 : _GEN_2391; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2456 = _T_177 ? _GEN_2184 : _GEN_2392; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2457 = _T_177 ? _GEN_2185 : _GEN_2393; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2458 = _T_177 ? _GEN_2186 : _GEN_2394; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2459 = _T_177 ? _GEN_2187 : _GEN_2395; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2460 = _T_177 ? _GEN_2188 : _GEN_2396; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2461 = _T_177 ? _GEN_2189 : _GEN_2397; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2462 = _T_177 ? _GEN_2190 : _GEN_2398; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2463 = _T_177 ? _GEN_2191 : _GEN_2399; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2464 = _T_177 ? _GEN_2192 : _GEN_2400; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2465 = _T_177 ? _GEN_2193 : _GEN_2401; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2466 = _T_177 ? _GEN_2194 : _GEN_2402; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2467 = _T_177 ? _GEN_2195 : _GEN_2403; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2468 = _T_177 ? _GEN_2196 : _GEN_2404; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2469 = _T_177 ? _GEN_2197 : _GEN_2405; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2470 = _T_177 ? _GEN_2198 : _GEN_2406; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2471 = _T_177 ? _GEN_2199 : _GEN_2407; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2472 = _T_177 ? _GEN_2200 : _GEN_2023; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2473 = _T_177 ? _GEN_2201 : _GEN_2024; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2474 = _T_177 ? _GEN_2202 : _GEN_2025; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2475 = _T_177 ? _GEN_2203 : _GEN_2026; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2476 = _T_177 ? _GEN_2204 : _GEN_2027; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2477 = _T_177 ? _GEN_2205 : _GEN_2028; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2478 = _T_177 ? _GEN_2206 : _GEN_2029; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2479 = _T_177 ? _GEN_2207 : _GEN_2030; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2480 = _T_177 ? _GEN_2208 : _GEN_2031; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2481 = _T_177 ? _GEN_2209 : _GEN_2032; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2482 = _T_177 ? _GEN_2210 : _GEN_2033; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2483 = _T_177 ? _GEN_2211 : _GEN_2034; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2484 = _T_177 ? _GEN_2212 : _GEN_2035; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2485 = _T_177 ? _GEN_2213 : _GEN_2036; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2486 = _T_177 ? _GEN_2214 : _GEN_2037; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2487 = _T_177 ? _GEN_2215 : _GEN_2038; // @[TBE.scala 114:59]
  wire  _T_287 = io_write_4_bits_command == 2'h1; // @[TBE.scala 136:44]
  wire  isAlloc_4 = _T_287 & io_write_4_valid; // @[TBE.scala 136:54]
  wire [31:0] _GEN_2489 = isAlloc_4 ? _GEN_2056 : _GEN_2424; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2490 = isAlloc_4 ? _GEN_2057 : _GEN_2425; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2491 = isAlloc_4 ? _GEN_2058 : _GEN_2426; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2492 = isAlloc_4 ? _GEN_2059 : _GEN_2427; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2493 = isAlloc_4 ? _GEN_2060 : _GEN_2428; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2494 = isAlloc_4 ? _GEN_2061 : _GEN_2429; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2495 = isAlloc_4 ? _GEN_2062 : _GEN_2430; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2496 = isAlloc_4 ? _GEN_2063 : _GEN_2431; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2497 = isAlloc_4 ? _GEN_2064 : _GEN_2432; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2498 = isAlloc_4 ? _GEN_2065 : _GEN_2433; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2499 = isAlloc_4 ? _GEN_2066 : _GEN_2434; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2500 = isAlloc_4 ? _GEN_2067 : _GEN_2435; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2501 = isAlloc_4 ? _GEN_2068 : _GEN_2436; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2502 = isAlloc_4 ? _GEN_2069 : _GEN_2437; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2503 = isAlloc_4 ? _GEN_2070 : _GEN_2438; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2504 = isAlloc_4 ? _GEN_2071 : _GEN_2439; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2505 = isAlloc_4 ? _GEN_2072 : _GEN_2440; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2506 = isAlloc_4 ? _GEN_2073 : _GEN_2441; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2507 = isAlloc_4 ? _GEN_2074 : _GEN_2442; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2508 = isAlloc_4 ? _GEN_2075 : _GEN_2443; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2509 = isAlloc_4 ? _GEN_2076 : _GEN_2444; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2510 = isAlloc_4 ? _GEN_2077 : _GEN_2445; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2511 = isAlloc_4 ? _GEN_2078 : _GEN_2446; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2512 = isAlloc_4 ? _GEN_2079 : _GEN_2447; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2513 = isAlloc_4 ? _GEN_2080 : _GEN_2448; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2514 = isAlloc_4 ? _GEN_2081 : _GEN_2449; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2515 = isAlloc_4 ? _GEN_2082 : _GEN_2450; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2516 = isAlloc_4 ? _GEN_2083 : _GEN_2451; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2517 = isAlloc_4 ? _GEN_2084 : _GEN_2452; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2518 = isAlloc_4 ? _GEN_2085 : _GEN_2453; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2519 = isAlloc_4 ? _GEN_2086 : _GEN_2454; // @[TBE.scala 109:24]
  wire [2:0] _GEN_2520 = isAlloc_4 ? _GEN_2087 : _GEN_2455; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2521 = isAlloc_4 ? _GEN_2088 : _GEN_2456; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2522 = isAlloc_4 ? _GEN_2089 : _GEN_2457; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2523 = isAlloc_4 ? _GEN_2090 : _GEN_2458; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2524 = isAlloc_4 ? _GEN_2091 : _GEN_2459; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2525 = isAlloc_4 ? _GEN_2092 : _GEN_2460; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2526 = isAlloc_4 ? _GEN_2093 : _GEN_2461; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2527 = isAlloc_4 ? _GEN_2094 : _GEN_2462; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2528 = isAlloc_4 ? _GEN_2095 : _GEN_2463; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2529 = isAlloc_4 ? _GEN_2096 : _GEN_2464; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2530 = isAlloc_4 ? _GEN_2097 : _GEN_2465; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2531 = isAlloc_4 ? _GEN_2098 : _GEN_2466; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2532 = isAlloc_4 ? _GEN_2099 : _GEN_2467; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2533 = isAlloc_4 ? _GEN_2100 : _GEN_2468; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2534 = isAlloc_4 ? _GEN_2101 : _GEN_2469; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2535 = isAlloc_4 ? _GEN_2102 : _GEN_2470; // @[TBE.scala 109:24]
  wire [1:0] _GEN_2536 = isAlloc_4 ? _GEN_2103 : _GEN_2471; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2537 = isAlloc_4 ? _GEN_2104 : _GEN_2472; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2538 = isAlloc_4 ? _GEN_2105 : _GEN_2473; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2539 = isAlloc_4 ? _GEN_2106 : _GEN_2474; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2540 = isAlloc_4 ? _GEN_2107 : _GEN_2475; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2541 = isAlloc_4 ? _GEN_2108 : _GEN_2476; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2542 = isAlloc_4 ? _GEN_2109 : _GEN_2477; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2543 = isAlloc_4 ? _GEN_2110 : _GEN_2478; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2544 = isAlloc_4 ? _GEN_2111 : _GEN_2479; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2545 = isAlloc_4 ? _GEN_2112 : _GEN_2480; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2546 = isAlloc_4 ? _GEN_2113 : _GEN_2481; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2547 = isAlloc_4 ? _GEN_2114 : _GEN_2482; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2548 = isAlloc_4 ? _GEN_2115 : _GEN_2483; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2549 = isAlloc_4 ? _GEN_2116 : _GEN_2484; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2550 = isAlloc_4 ? _GEN_2117 : _GEN_2485; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2551 = isAlloc_4 ? _GEN_2118 : _GEN_2486; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2552 = isAlloc_4 ? _GEN_2119 : _GEN_2487; // @[TBE.scala 109:24]
  wire  _GEN_2553 = isAlloc_4 ? _GEN_2120 : _GEN_2408; // @[TBE.scala 109:24]
  wire  _GEN_2554 = isAlloc_4 ? _GEN_2121 : _GEN_2409; // @[TBE.scala 109:24]
  wire  _GEN_2555 = isAlloc_4 ? _GEN_2122 : _GEN_2410; // @[TBE.scala 109:24]
  wire  _GEN_2556 = isAlloc_4 ? _GEN_2123 : _GEN_2411; // @[TBE.scala 109:24]
  wire  _GEN_2557 = isAlloc_4 ? _GEN_2124 : _GEN_2412; // @[TBE.scala 109:24]
  wire  _GEN_2558 = isAlloc_4 ? _GEN_2125 : _GEN_2413; // @[TBE.scala 109:24]
  wire  _GEN_2559 = isAlloc_4 ? _GEN_2126 : _GEN_2414; // @[TBE.scala 109:24]
  wire  _GEN_2560 = isAlloc_4 ? _GEN_2127 : _GEN_2415; // @[TBE.scala 109:24]
  wire  _GEN_2561 = isAlloc_4 ? _GEN_2128 : _GEN_2416; // @[TBE.scala 109:24]
  wire  _GEN_2562 = isAlloc_4 ? _GEN_2129 : _GEN_2417; // @[TBE.scala 109:24]
  wire  _GEN_2563 = isAlloc_4 ? _GEN_2130 : _GEN_2418; // @[TBE.scala 109:24]
  wire  _GEN_2564 = isAlloc_4 ? _GEN_2131 : _GEN_2419; // @[TBE.scala 109:24]
  wire  _GEN_2565 = isAlloc_4 ? _GEN_2132 : _GEN_2420; // @[TBE.scala 109:24]
  wire  _GEN_2566 = isAlloc_4 ? _GEN_2133 : _GEN_2421; // @[TBE.scala 109:24]
  wire  _GEN_2567 = isAlloc_4 ? _GEN_2134 : _GEN_2422; // @[TBE.scala 109:24]
  wire  _GEN_2568 = isAlloc_4 ? _GEN_2135 : _GEN_2423; // @[TBE.scala 109:24]
  wire [31:0] _GEN_2570 = 4'h0 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2489; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2571 = 4'h1 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2490; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2572 = 4'h2 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2491; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2573 = 4'h3 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2492; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2574 = 4'h4 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2493; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2575 = 4'h5 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2494; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2576 = 4'h6 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2495; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2577 = 4'h7 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2496; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2578 = 4'h8 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2497; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2579 = 4'h9 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2498; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2580 = 4'ha == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2499; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2581 = 4'hb == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2500; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2582 = 4'hc == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2501; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2583 = 4'hd == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2502; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2584 = 4'he == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2503; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2585 = 4'hf == idxAlloc[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2504; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2586 = 4'h0 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2505; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2587 = 4'h1 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2506; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2588 = 4'h2 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2507; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2589 = 4'h3 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2508; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2590 = 4'h4 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2509; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2591 = 4'h5 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2510; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2592 = 4'h6 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2511; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2593 = 4'h7 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2512; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2594 = 4'h8 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2513; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2595 = 4'h9 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2514; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2596 = 4'ha == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2515; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2597 = 4'hb == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2516; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2598 = 4'hc == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2517; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2599 = 4'hd == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2518; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2600 = 4'he == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2519; // @[TBE.scala 110:27]
  wire [2:0] _GEN_2601 = 4'hf == idxAlloc[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2520; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2602 = 4'h0 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2521; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2603 = 4'h1 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2522; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2604 = 4'h2 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2523; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2605 = 4'h3 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2524; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2606 = 4'h4 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2525; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2607 = 4'h5 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2526; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2608 = 4'h6 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2527; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2609 = 4'h7 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2528; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2610 = 4'h8 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2529; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2611 = 4'h9 == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2530; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2612 = 4'ha == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2531; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2613 = 4'hb == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2532; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2614 = 4'hc == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2533; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2615 = 4'hd == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2534; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2616 = 4'he == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2535; // @[TBE.scala 110:27]
  wire [1:0] _GEN_2617 = 4'hf == idxAlloc[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2536; // @[TBE.scala 110:27]
  wire [31:0] _GEN_2618 = 4'h0 == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2537; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2619 = 4'h1 == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2538; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2620 = 4'h2 == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2539; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2621 = 4'h3 == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2540; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2622 = 4'h4 == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2541; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2623 = 4'h5 == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2542; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2624 = 4'h6 == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2543; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2625 = 4'h7 == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2544; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2626 = 4'h8 == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2545; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2627 = 4'h9 == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2546; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2628 = 4'ha == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2547; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2629 = 4'hb == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2548; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2630 = 4'hc == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2549; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2631 = 4'hd == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2550; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2632 = 4'he == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2551; // @[TBE.scala 111:25]
  wire [31:0] _GEN_2633 = 4'hf == idxAlloc[3:0] ? io_write_5_bits_addr[31:0] : _GEN_2552; // @[TBE.scala 111:25]
  wire  _GEN_2634 = _GEN_4161 | _GEN_2553; // @[TBE.scala 112:26]
  wire  _GEN_2635 = _GEN_4162 | _GEN_2554; // @[TBE.scala 112:26]
  wire  _GEN_2636 = _GEN_4163 | _GEN_2555; // @[TBE.scala 112:26]
  wire  _GEN_2637 = _GEN_4164 | _GEN_2556; // @[TBE.scala 112:26]
  wire  _GEN_2638 = _GEN_4165 | _GEN_2557; // @[TBE.scala 112:26]
  wire  _GEN_2639 = _GEN_4166 | _GEN_2558; // @[TBE.scala 112:26]
  wire  _GEN_2640 = _GEN_4167 | _GEN_2559; // @[TBE.scala 112:26]
  wire  _GEN_2641 = _GEN_4168 | _GEN_2560; // @[TBE.scala 112:26]
  wire  _GEN_2642 = _GEN_4169 | _GEN_2561; // @[TBE.scala 112:26]
  wire  _GEN_2643 = _GEN_4170 | _GEN_2562; // @[TBE.scala 112:26]
  wire  _GEN_2644 = _GEN_4171 | _GEN_2563; // @[TBE.scala 112:26]
  wire  _GEN_2645 = _GEN_4172 | _GEN_2564; // @[TBE.scala 112:26]
  wire  _GEN_2646 = _GEN_4173 | _GEN_2565; // @[TBE.scala 112:26]
  wire  _GEN_2647 = _GEN_4174 | _GEN_2566; // @[TBE.scala 112:26]
  wire  _GEN_2648 = _GEN_4175 | _GEN_2567; // @[TBE.scala 112:26]
  wire  _GEN_2649 = _GEN_4176 | _GEN_2568; // @[TBE.scala 112:26]
  wire  _T_295 = io_write_5_bits_command == 2'h2; // @[TBE.scala 137:46]
  wire  isDealloc_5 = _T_295 & io_write_5_valid; // @[TBE.scala 137:58]
  wire  _T_199 = isDealloc_5 & finder_5_io_value_valid; // @[TBE.scala 114:31]
  wire [4:0] idxUpdate_5 = {{1'd0}, finder_5_io_value_bits}; // @[TBE.scala 73:23 TBE.scala 104:18]
  wire  _GEN_2650 = 4'h0 == idxUpdate_5[3:0] ? 1'h0 : _GEN_2553; // @[TBE.scala 115:30]
  wire  _GEN_2651 = 4'h1 == idxUpdate_5[3:0] ? 1'h0 : _GEN_2554; // @[TBE.scala 115:30]
  wire  _GEN_2652 = 4'h2 == idxUpdate_5[3:0] ? 1'h0 : _GEN_2555; // @[TBE.scala 115:30]
  wire  _GEN_2653 = 4'h3 == idxUpdate_5[3:0] ? 1'h0 : _GEN_2556; // @[TBE.scala 115:30]
  wire  _GEN_2654 = 4'h4 == idxUpdate_5[3:0] ? 1'h0 : _GEN_2557; // @[TBE.scala 115:30]
  wire  _GEN_2655 = 4'h5 == idxUpdate_5[3:0] ? 1'h0 : _GEN_2558; // @[TBE.scala 115:30]
  wire  _GEN_2656 = 4'h6 == idxUpdate_5[3:0] ? 1'h0 : _GEN_2559; // @[TBE.scala 115:30]
  wire  _GEN_2657 = 4'h7 == idxUpdate_5[3:0] ? 1'h0 : _GEN_2560; // @[TBE.scala 115:30]
  wire  _GEN_2658 = 4'h8 == idxUpdate_5[3:0] ? 1'h0 : _GEN_2561; // @[TBE.scala 115:30]
  wire  _GEN_2659 = 4'h9 == idxUpdate_5[3:0] ? 1'h0 : _GEN_2562; // @[TBE.scala 115:30]
  wire  _GEN_2660 = 4'ha == idxUpdate_5[3:0] ? 1'h0 : _GEN_2563; // @[TBE.scala 115:30]
  wire  _GEN_2661 = 4'hb == idxUpdate_5[3:0] ? 1'h0 : _GEN_2564; // @[TBE.scala 115:30]
  wire  _GEN_2662 = 4'hc == idxUpdate_5[3:0] ? 1'h0 : _GEN_2565; // @[TBE.scala 115:30]
  wire  _GEN_2663 = 4'hd == idxUpdate_5[3:0] ? 1'h0 : _GEN_2566; // @[TBE.scala 115:30]
  wire  _GEN_2664 = 4'he == idxUpdate_5[3:0] ? 1'h0 : _GEN_2567; // @[TBE.scala 115:30]
  wire  _GEN_2665 = 4'hf == idxUpdate_5[3:0] ? 1'h0 : _GEN_2568; // @[TBE.scala 115:30]
  wire [31:0] _GEN_2666 = 4'h0 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2489; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2667 = 4'h1 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2490; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2668 = 4'h2 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2491; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2669 = 4'h3 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2492; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2670 = 4'h4 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2493; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2671 = 4'h5 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2494; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2672 = 4'h6 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2495; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2673 = 4'h7 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2496; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2674 = 4'h8 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2497; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2675 = 4'h9 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2498; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2676 = 4'ha == idxUpdate_5[3:0] ? 32'h0 : _GEN_2499; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2677 = 4'hb == idxUpdate_5[3:0] ? 32'h0 : _GEN_2500; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2678 = 4'hc == idxUpdate_5[3:0] ? 32'h0 : _GEN_2501; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2679 = 4'hd == idxUpdate_5[3:0] ? 32'h0 : _GEN_2502; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2680 = 4'he == idxUpdate_5[3:0] ? 32'h0 : _GEN_2503; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2681 = 4'hf == idxUpdate_5[3:0] ? 32'h0 : _GEN_2504; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2682 = 4'h0 == idxUpdate_5[3:0] ? 3'h2 : _GEN_2505; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2683 = 4'h1 == idxUpdate_5[3:0] ? 3'h2 : _GEN_2506; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2684 = 4'h2 == idxUpdate_5[3:0] ? 3'h2 : _GEN_2507; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2685 = 4'h3 == idxUpdate_5[3:0] ? 3'h2 : _GEN_2508; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2686 = 4'h4 == idxUpdate_5[3:0] ? 3'h2 : _GEN_2509; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2687 = 4'h5 == idxUpdate_5[3:0] ? 3'h2 : _GEN_2510; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2688 = 4'h6 == idxUpdate_5[3:0] ? 3'h2 : _GEN_2511; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2689 = 4'h7 == idxUpdate_5[3:0] ? 3'h2 : _GEN_2512; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2690 = 4'h8 == idxUpdate_5[3:0] ? 3'h2 : _GEN_2513; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2691 = 4'h9 == idxUpdate_5[3:0] ? 3'h2 : _GEN_2514; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2692 = 4'ha == idxUpdate_5[3:0] ? 3'h2 : _GEN_2515; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2693 = 4'hb == idxUpdate_5[3:0] ? 3'h2 : _GEN_2516; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2694 = 4'hc == idxUpdate_5[3:0] ? 3'h2 : _GEN_2517; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2695 = 4'hd == idxUpdate_5[3:0] ? 3'h2 : _GEN_2518; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2696 = 4'he == idxUpdate_5[3:0] ? 3'h2 : _GEN_2519; // @[TBE.scala 116:31]
  wire [2:0] _GEN_2697 = 4'hf == idxUpdate_5[3:0] ? 3'h2 : _GEN_2520; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2698 = 4'h0 == idxUpdate_5[3:0] ? 2'h0 : _GEN_2521; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2699 = 4'h1 == idxUpdate_5[3:0] ? 2'h0 : _GEN_2522; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2700 = 4'h2 == idxUpdate_5[3:0] ? 2'h0 : _GEN_2523; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2701 = 4'h3 == idxUpdate_5[3:0] ? 2'h0 : _GEN_2524; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2702 = 4'h4 == idxUpdate_5[3:0] ? 2'h0 : _GEN_2525; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2703 = 4'h5 == idxUpdate_5[3:0] ? 2'h0 : _GEN_2526; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2704 = 4'h6 == idxUpdate_5[3:0] ? 2'h0 : _GEN_2527; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2705 = 4'h7 == idxUpdate_5[3:0] ? 2'h0 : _GEN_2528; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2706 = 4'h8 == idxUpdate_5[3:0] ? 2'h0 : _GEN_2529; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2707 = 4'h9 == idxUpdate_5[3:0] ? 2'h0 : _GEN_2530; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2708 = 4'ha == idxUpdate_5[3:0] ? 2'h0 : _GEN_2531; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2709 = 4'hb == idxUpdate_5[3:0] ? 2'h0 : _GEN_2532; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2710 = 4'hc == idxUpdate_5[3:0] ? 2'h0 : _GEN_2533; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2711 = 4'hd == idxUpdate_5[3:0] ? 2'h0 : _GEN_2534; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2712 = 4'he == idxUpdate_5[3:0] ? 2'h0 : _GEN_2535; // @[TBE.scala 116:31]
  wire [1:0] _GEN_2713 = 4'hf == idxUpdate_5[3:0] ? 2'h0 : _GEN_2536; // @[TBE.scala 116:31]
  wire [31:0] _GEN_2714 = 4'h0 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2537; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2715 = 4'h1 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2538; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2716 = 4'h2 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2539; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2717 = 4'h3 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2540; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2718 = 4'h4 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2541; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2719 = 4'h5 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2542; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2720 = 4'h6 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2543; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2721 = 4'h7 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2544; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2722 = 4'h8 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2545; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2723 = 4'h9 == idxUpdate_5[3:0] ? 32'h0 : _GEN_2546; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2724 = 4'ha == idxUpdate_5[3:0] ? 32'h0 : _GEN_2547; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2725 = 4'hb == idxUpdate_5[3:0] ? 32'h0 : _GEN_2548; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2726 = 4'hc == idxUpdate_5[3:0] ? 32'h0 : _GEN_2549; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2727 = 4'hd == idxUpdate_5[3:0] ? 32'h0 : _GEN_2550; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2728 = 4'he == idxUpdate_5[3:0] ? 32'h0 : _GEN_2551; // @[TBE.scala 117:29]
  wire [31:0] _GEN_2729 = 4'hf == idxUpdate_5[3:0] ? 32'h0 : _GEN_2552; // @[TBE.scala 117:29]
  wire  _T_297 = io_write_5_bits_command == 2'h3; // @[TBE.scala 138:44]
  wire  isWrite_5 = _T_297 & io_write_5_valid; // @[TBE.scala 138:55]
  wire  _T_207 = isWrite_5 & finder_5_io_value_valid; // @[TBE.scala 119:29]
  wire  _T_208 = ~io_write_5_bits_mask; // @[TBE.scala 120:35]
  wire [31:0] _GEN_2730 = 4'h0 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2489; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2731 = 4'h1 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2490; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2732 = 4'h2 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2491; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2733 = 4'h3 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2492; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2734 = 4'h4 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2493; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2735 = 4'h5 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2494; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2736 = 4'h6 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2495; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2737 = 4'h7 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2496; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2738 = 4'h8 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2497; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2739 = 4'h9 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2498; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2740 = 4'ha == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2499; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2741 = 4'hb == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2500; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2742 = 4'hc == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2501; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2743 = 4'hd == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2502; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2744 = 4'he == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2503; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2745 = 4'hf == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_fields_0 : _GEN_2504; // @[TBE.scala 121:63]
  wire [31:0] _GEN_2751 = 4'h1 == idxUpdate_5[3:0] ? TBEMemory_1_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2754 = 4'h2 == idxUpdate_5[3:0] ? TBEMemory_2_fields_0 : _GEN_2751; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2757 = 4'h3 == idxUpdate_5[3:0] ? TBEMemory_3_fields_0 : _GEN_2754; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2760 = 4'h4 == idxUpdate_5[3:0] ? TBEMemory_4_fields_0 : _GEN_2757; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2763 = 4'h5 == idxUpdate_5[3:0] ? TBEMemory_5_fields_0 : _GEN_2760; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2766 = 4'h6 == idxUpdate_5[3:0] ? TBEMemory_6_fields_0 : _GEN_2763; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2769 = 4'h7 == idxUpdate_5[3:0] ? TBEMemory_7_fields_0 : _GEN_2766; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2772 = 4'h8 == idxUpdate_5[3:0] ? TBEMemory_8_fields_0 : _GEN_2769; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2775 = 4'h9 == idxUpdate_5[3:0] ? TBEMemory_9_fields_0 : _GEN_2772; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2778 = 4'ha == idxUpdate_5[3:0] ? TBEMemory_10_fields_0 : _GEN_2775; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2781 = 4'hb == idxUpdate_5[3:0] ? TBEMemory_11_fields_0 : _GEN_2778; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2784 = 4'hc == idxUpdate_5[3:0] ? TBEMemory_12_fields_0 : _GEN_2781; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2787 = 4'hd == idxUpdate_5[3:0] ? TBEMemory_13_fields_0 : _GEN_2784; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2790 = 4'he == idxUpdate_5[3:0] ? TBEMemory_14_fields_0 : _GEN_2787; // @[TBE.scala 122:15]
  wire [31:0] _GEN_2793 = 4'hf == idxUpdate_5[3:0] ? TBEMemory_15_fields_0 : _GEN_2790; // @[TBE.scala 122:15]
  wire [2:0] _GEN_2794 = 4'h0 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2505; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2795 = 4'h1 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2506; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2796 = 4'h2 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2507; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2797 = 4'h3 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2508; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2798 = 4'h4 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2509; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2799 = 4'h5 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2510; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2800 = 4'h6 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2511; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2801 = 4'h7 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2512; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2802 = 4'h8 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2513; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2803 = 4'h9 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2514; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2804 = 4'ha == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2515; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2805 = 4'hb == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2516; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2806 = 4'hc == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2517; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2807 = 4'hd == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2518; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2808 = 4'he == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2519; // @[TBE.scala 124:37]
  wire [2:0] _GEN_2809 = 4'hf == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_way : _GEN_2520; // @[TBE.scala 124:37]
  wire [1:0] _GEN_2810 = 4'h0 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2521; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2811 = 4'h1 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2522; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2812 = 4'h2 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2523; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2813 = 4'h3 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2524; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2814 = 4'h4 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2525; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2815 = 4'h5 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2526; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2816 = 4'h6 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2527; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2817 = 4'h7 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2528; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2818 = 4'h8 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2529; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2819 = 4'h9 == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2530; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2820 = 4'ha == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2531; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2821 = 4'hb == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2532; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2822 = 4'hc == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2533; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2823 = 4'hd == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2534; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2824 = 4'he == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2535; // @[TBE.scala 125:39]
  wire [1:0] _GEN_2825 = 4'hf == idxUpdate_5[3:0] ? io_write_5_bits_inputTBE_state_state : _GEN_2536; // @[TBE.scala 125:39]
  wire [31:0] _GEN_2826 = _T_208 ? _GEN_2730 : _GEN_2489; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2827 = _T_208 ? _GEN_2731 : _GEN_2490; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2828 = _T_208 ? _GEN_2732 : _GEN_2491; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2829 = _T_208 ? _GEN_2733 : _GEN_2492; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2830 = _T_208 ? _GEN_2734 : _GEN_2493; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2831 = _T_208 ? _GEN_2735 : _GEN_2494; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2832 = _T_208 ? _GEN_2736 : _GEN_2495; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2833 = _T_208 ? _GEN_2737 : _GEN_2496; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2834 = _T_208 ? _GEN_2738 : _GEN_2497; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2835 = _T_208 ? _GEN_2739 : _GEN_2498; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2836 = _T_208 ? _GEN_2740 : _GEN_2499; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2837 = _T_208 ? _GEN_2741 : _GEN_2500; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2838 = _T_208 ? _GEN_2742 : _GEN_2501; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2839 = _T_208 ? _GEN_2743 : _GEN_2502; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2840 = _T_208 ? _GEN_2744 : _GEN_2503; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2841 = _T_208 ? _GEN_2745 : _GEN_2504; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2842 = _T_208 ? _GEN_2505 : _GEN_2794; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2843 = _T_208 ? _GEN_2506 : _GEN_2795; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2844 = _T_208 ? _GEN_2507 : _GEN_2796; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2845 = _T_208 ? _GEN_2508 : _GEN_2797; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2846 = _T_208 ? _GEN_2509 : _GEN_2798; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2847 = _T_208 ? _GEN_2510 : _GEN_2799; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2848 = _T_208 ? _GEN_2511 : _GEN_2800; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2849 = _T_208 ? _GEN_2512 : _GEN_2801; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2850 = _T_208 ? _GEN_2513 : _GEN_2802; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2851 = _T_208 ? _GEN_2514 : _GEN_2803; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2852 = _T_208 ? _GEN_2515 : _GEN_2804; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2853 = _T_208 ? _GEN_2516 : _GEN_2805; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2854 = _T_208 ? _GEN_2517 : _GEN_2806; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2855 = _T_208 ? _GEN_2518 : _GEN_2807; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2856 = _T_208 ? _GEN_2519 : _GEN_2808; // @[TBE.scala 120:53]
  wire [2:0] _GEN_2857 = _T_208 ? _GEN_2520 : _GEN_2809; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2858 = _T_208 ? _GEN_2521 : _GEN_2810; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2859 = _T_208 ? _GEN_2522 : _GEN_2811; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2860 = _T_208 ? _GEN_2523 : _GEN_2812; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2861 = _T_208 ? _GEN_2524 : _GEN_2813; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2862 = _T_208 ? _GEN_2525 : _GEN_2814; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2863 = _T_208 ? _GEN_2526 : _GEN_2815; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2864 = _T_208 ? _GEN_2527 : _GEN_2816; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2865 = _T_208 ? _GEN_2528 : _GEN_2817; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2866 = _T_208 ? _GEN_2529 : _GEN_2818; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2867 = _T_208 ? _GEN_2530 : _GEN_2819; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2868 = _T_208 ? _GEN_2531 : _GEN_2820; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2869 = _T_208 ? _GEN_2532 : _GEN_2821; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2870 = _T_208 ? _GEN_2533 : _GEN_2822; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2871 = _T_208 ? _GEN_2534 : _GEN_2823; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2872 = _T_208 ? _GEN_2535 : _GEN_2824; // @[TBE.scala 120:53]
  wire [1:0] _GEN_2873 = _T_208 ? _GEN_2536 : _GEN_2825; // @[TBE.scala 120:53]
  wire [31:0] _GEN_2874 = _T_207 ? _GEN_2826 : _GEN_2489; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2875 = _T_207 ? _GEN_2827 : _GEN_2490; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2876 = _T_207 ? _GEN_2828 : _GEN_2491; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2877 = _T_207 ? _GEN_2829 : _GEN_2492; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2878 = _T_207 ? _GEN_2830 : _GEN_2493; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2879 = _T_207 ? _GEN_2831 : _GEN_2494; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2880 = _T_207 ? _GEN_2832 : _GEN_2495; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2881 = _T_207 ? _GEN_2833 : _GEN_2496; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2882 = _T_207 ? _GEN_2834 : _GEN_2497; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2883 = _T_207 ? _GEN_2835 : _GEN_2498; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2884 = _T_207 ? _GEN_2836 : _GEN_2499; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2885 = _T_207 ? _GEN_2837 : _GEN_2500; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2886 = _T_207 ? _GEN_2838 : _GEN_2501; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2887 = _T_207 ? _GEN_2839 : _GEN_2502; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2888 = _T_207 ? _GEN_2840 : _GEN_2503; // @[TBE.scala 119:57]
  wire [31:0] _GEN_2889 = _T_207 ? _GEN_2841 : _GEN_2504; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2890 = _T_207 ? _GEN_2842 : _GEN_2505; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2891 = _T_207 ? _GEN_2843 : _GEN_2506; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2892 = _T_207 ? _GEN_2844 : _GEN_2507; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2893 = _T_207 ? _GEN_2845 : _GEN_2508; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2894 = _T_207 ? _GEN_2846 : _GEN_2509; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2895 = _T_207 ? _GEN_2847 : _GEN_2510; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2896 = _T_207 ? _GEN_2848 : _GEN_2511; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2897 = _T_207 ? _GEN_2849 : _GEN_2512; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2898 = _T_207 ? _GEN_2850 : _GEN_2513; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2899 = _T_207 ? _GEN_2851 : _GEN_2514; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2900 = _T_207 ? _GEN_2852 : _GEN_2515; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2901 = _T_207 ? _GEN_2853 : _GEN_2516; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2902 = _T_207 ? _GEN_2854 : _GEN_2517; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2903 = _T_207 ? _GEN_2855 : _GEN_2518; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2904 = _T_207 ? _GEN_2856 : _GEN_2519; // @[TBE.scala 119:57]
  wire [2:0] _GEN_2905 = _T_207 ? _GEN_2857 : _GEN_2520; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2906 = _T_207 ? _GEN_2858 : _GEN_2521; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2907 = _T_207 ? _GEN_2859 : _GEN_2522; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2908 = _T_207 ? _GEN_2860 : _GEN_2523; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2909 = _T_207 ? _GEN_2861 : _GEN_2524; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2910 = _T_207 ? _GEN_2862 : _GEN_2525; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2911 = _T_207 ? _GEN_2863 : _GEN_2526; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2912 = _T_207 ? _GEN_2864 : _GEN_2527; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2913 = _T_207 ? _GEN_2865 : _GEN_2528; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2914 = _T_207 ? _GEN_2866 : _GEN_2529; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2915 = _T_207 ? _GEN_2867 : _GEN_2530; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2916 = _T_207 ? _GEN_2868 : _GEN_2531; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2917 = _T_207 ? _GEN_2869 : _GEN_2532; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2918 = _T_207 ? _GEN_2870 : _GEN_2533; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2919 = _T_207 ? _GEN_2871 : _GEN_2534; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2920 = _T_207 ? _GEN_2872 : _GEN_2535; // @[TBE.scala 119:57]
  wire [1:0] _GEN_2921 = _T_207 ? _GEN_2873 : _GEN_2536; // @[TBE.scala 119:57]
  wire  _GEN_2922 = _T_199 ? _GEN_2650 : _GEN_2553; // @[TBE.scala 114:59]
  wire  _GEN_2923 = _T_199 ? _GEN_2651 : _GEN_2554; // @[TBE.scala 114:59]
  wire  _GEN_2924 = _T_199 ? _GEN_2652 : _GEN_2555; // @[TBE.scala 114:59]
  wire  _GEN_2925 = _T_199 ? _GEN_2653 : _GEN_2556; // @[TBE.scala 114:59]
  wire  _GEN_2926 = _T_199 ? _GEN_2654 : _GEN_2557; // @[TBE.scala 114:59]
  wire  _GEN_2927 = _T_199 ? _GEN_2655 : _GEN_2558; // @[TBE.scala 114:59]
  wire  _GEN_2928 = _T_199 ? _GEN_2656 : _GEN_2559; // @[TBE.scala 114:59]
  wire  _GEN_2929 = _T_199 ? _GEN_2657 : _GEN_2560; // @[TBE.scala 114:59]
  wire  _GEN_2930 = _T_199 ? _GEN_2658 : _GEN_2561; // @[TBE.scala 114:59]
  wire  _GEN_2931 = _T_199 ? _GEN_2659 : _GEN_2562; // @[TBE.scala 114:59]
  wire  _GEN_2932 = _T_199 ? _GEN_2660 : _GEN_2563; // @[TBE.scala 114:59]
  wire  _GEN_2933 = _T_199 ? _GEN_2661 : _GEN_2564; // @[TBE.scala 114:59]
  wire  _GEN_2934 = _T_199 ? _GEN_2662 : _GEN_2565; // @[TBE.scala 114:59]
  wire  _GEN_2935 = _T_199 ? _GEN_2663 : _GEN_2566; // @[TBE.scala 114:59]
  wire  _GEN_2936 = _T_199 ? _GEN_2664 : _GEN_2567; // @[TBE.scala 114:59]
  wire  _GEN_2937 = _T_199 ? _GEN_2665 : _GEN_2568; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2938 = _T_199 ? _GEN_2666 : _GEN_2874; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2939 = _T_199 ? _GEN_2667 : _GEN_2875; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2940 = _T_199 ? _GEN_2668 : _GEN_2876; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2941 = _T_199 ? _GEN_2669 : _GEN_2877; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2942 = _T_199 ? _GEN_2670 : _GEN_2878; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2943 = _T_199 ? _GEN_2671 : _GEN_2879; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2944 = _T_199 ? _GEN_2672 : _GEN_2880; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2945 = _T_199 ? _GEN_2673 : _GEN_2881; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2946 = _T_199 ? _GEN_2674 : _GEN_2882; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2947 = _T_199 ? _GEN_2675 : _GEN_2883; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2948 = _T_199 ? _GEN_2676 : _GEN_2884; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2949 = _T_199 ? _GEN_2677 : _GEN_2885; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2950 = _T_199 ? _GEN_2678 : _GEN_2886; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2951 = _T_199 ? _GEN_2679 : _GEN_2887; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2952 = _T_199 ? _GEN_2680 : _GEN_2888; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2953 = _T_199 ? _GEN_2681 : _GEN_2889; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2954 = _T_199 ? _GEN_2682 : _GEN_2890; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2955 = _T_199 ? _GEN_2683 : _GEN_2891; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2956 = _T_199 ? _GEN_2684 : _GEN_2892; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2957 = _T_199 ? _GEN_2685 : _GEN_2893; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2958 = _T_199 ? _GEN_2686 : _GEN_2894; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2959 = _T_199 ? _GEN_2687 : _GEN_2895; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2960 = _T_199 ? _GEN_2688 : _GEN_2896; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2961 = _T_199 ? _GEN_2689 : _GEN_2897; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2962 = _T_199 ? _GEN_2690 : _GEN_2898; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2963 = _T_199 ? _GEN_2691 : _GEN_2899; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2964 = _T_199 ? _GEN_2692 : _GEN_2900; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2965 = _T_199 ? _GEN_2693 : _GEN_2901; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2966 = _T_199 ? _GEN_2694 : _GEN_2902; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2967 = _T_199 ? _GEN_2695 : _GEN_2903; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2968 = _T_199 ? _GEN_2696 : _GEN_2904; // @[TBE.scala 114:59]
  wire [2:0] _GEN_2969 = _T_199 ? _GEN_2697 : _GEN_2905; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2970 = _T_199 ? _GEN_2698 : _GEN_2906; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2971 = _T_199 ? _GEN_2699 : _GEN_2907; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2972 = _T_199 ? _GEN_2700 : _GEN_2908; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2973 = _T_199 ? _GEN_2701 : _GEN_2909; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2974 = _T_199 ? _GEN_2702 : _GEN_2910; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2975 = _T_199 ? _GEN_2703 : _GEN_2911; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2976 = _T_199 ? _GEN_2704 : _GEN_2912; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2977 = _T_199 ? _GEN_2705 : _GEN_2913; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2978 = _T_199 ? _GEN_2706 : _GEN_2914; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2979 = _T_199 ? _GEN_2707 : _GEN_2915; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2980 = _T_199 ? _GEN_2708 : _GEN_2916; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2981 = _T_199 ? _GEN_2709 : _GEN_2917; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2982 = _T_199 ? _GEN_2710 : _GEN_2918; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2983 = _T_199 ? _GEN_2711 : _GEN_2919; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2984 = _T_199 ? _GEN_2712 : _GEN_2920; // @[TBE.scala 114:59]
  wire [1:0] _GEN_2985 = _T_199 ? _GEN_2713 : _GEN_2921; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2986 = _T_199 ? _GEN_2714 : _GEN_2537; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2987 = _T_199 ? _GEN_2715 : _GEN_2538; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2988 = _T_199 ? _GEN_2716 : _GEN_2539; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2989 = _T_199 ? _GEN_2717 : _GEN_2540; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2990 = _T_199 ? _GEN_2718 : _GEN_2541; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2991 = _T_199 ? _GEN_2719 : _GEN_2542; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2992 = _T_199 ? _GEN_2720 : _GEN_2543; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2993 = _T_199 ? _GEN_2721 : _GEN_2544; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2994 = _T_199 ? _GEN_2722 : _GEN_2545; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2995 = _T_199 ? _GEN_2723 : _GEN_2546; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2996 = _T_199 ? _GEN_2724 : _GEN_2547; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2997 = _T_199 ? _GEN_2725 : _GEN_2548; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2998 = _T_199 ? _GEN_2726 : _GEN_2549; // @[TBE.scala 114:59]
  wire [31:0] _GEN_2999 = _T_199 ? _GEN_2727 : _GEN_2550; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3000 = _T_199 ? _GEN_2728 : _GEN_2551; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3001 = _T_199 ? _GEN_2729 : _GEN_2552; // @[TBE.scala 114:59]
  wire  _T_293 = io_write_5_bits_command == 2'h1; // @[TBE.scala 136:44]
  wire  isAlloc_5 = _T_293 & io_write_5_valid; // @[TBE.scala 136:54]
  wire [31:0] _GEN_3003 = isAlloc_5 ? _GEN_2570 : _GEN_2938; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3004 = isAlloc_5 ? _GEN_2571 : _GEN_2939; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3005 = isAlloc_5 ? _GEN_2572 : _GEN_2940; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3006 = isAlloc_5 ? _GEN_2573 : _GEN_2941; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3007 = isAlloc_5 ? _GEN_2574 : _GEN_2942; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3008 = isAlloc_5 ? _GEN_2575 : _GEN_2943; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3009 = isAlloc_5 ? _GEN_2576 : _GEN_2944; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3010 = isAlloc_5 ? _GEN_2577 : _GEN_2945; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3011 = isAlloc_5 ? _GEN_2578 : _GEN_2946; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3012 = isAlloc_5 ? _GEN_2579 : _GEN_2947; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3013 = isAlloc_5 ? _GEN_2580 : _GEN_2948; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3014 = isAlloc_5 ? _GEN_2581 : _GEN_2949; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3015 = isAlloc_5 ? _GEN_2582 : _GEN_2950; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3016 = isAlloc_5 ? _GEN_2583 : _GEN_2951; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3017 = isAlloc_5 ? _GEN_2584 : _GEN_2952; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3018 = isAlloc_5 ? _GEN_2585 : _GEN_2953; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3019 = isAlloc_5 ? _GEN_2586 : _GEN_2954; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3020 = isAlloc_5 ? _GEN_2587 : _GEN_2955; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3021 = isAlloc_5 ? _GEN_2588 : _GEN_2956; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3022 = isAlloc_5 ? _GEN_2589 : _GEN_2957; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3023 = isAlloc_5 ? _GEN_2590 : _GEN_2958; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3024 = isAlloc_5 ? _GEN_2591 : _GEN_2959; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3025 = isAlloc_5 ? _GEN_2592 : _GEN_2960; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3026 = isAlloc_5 ? _GEN_2593 : _GEN_2961; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3027 = isAlloc_5 ? _GEN_2594 : _GEN_2962; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3028 = isAlloc_5 ? _GEN_2595 : _GEN_2963; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3029 = isAlloc_5 ? _GEN_2596 : _GEN_2964; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3030 = isAlloc_5 ? _GEN_2597 : _GEN_2965; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3031 = isAlloc_5 ? _GEN_2598 : _GEN_2966; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3032 = isAlloc_5 ? _GEN_2599 : _GEN_2967; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3033 = isAlloc_5 ? _GEN_2600 : _GEN_2968; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3034 = isAlloc_5 ? _GEN_2601 : _GEN_2969; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3035 = isAlloc_5 ? _GEN_2602 : _GEN_2970; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3036 = isAlloc_5 ? _GEN_2603 : _GEN_2971; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3037 = isAlloc_5 ? _GEN_2604 : _GEN_2972; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3038 = isAlloc_5 ? _GEN_2605 : _GEN_2973; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3039 = isAlloc_5 ? _GEN_2606 : _GEN_2974; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3040 = isAlloc_5 ? _GEN_2607 : _GEN_2975; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3041 = isAlloc_5 ? _GEN_2608 : _GEN_2976; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3042 = isAlloc_5 ? _GEN_2609 : _GEN_2977; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3043 = isAlloc_5 ? _GEN_2610 : _GEN_2978; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3044 = isAlloc_5 ? _GEN_2611 : _GEN_2979; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3045 = isAlloc_5 ? _GEN_2612 : _GEN_2980; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3046 = isAlloc_5 ? _GEN_2613 : _GEN_2981; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3047 = isAlloc_5 ? _GEN_2614 : _GEN_2982; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3048 = isAlloc_5 ? _GEN_2615 : _GEN_2983; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3049 = isAlloc_5 ? _GEN_2616 : _GEN_2984; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3050 = isAlloc_5 ? _GEN_2617 : _GEN_2985; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3051 = isAlloc_5 ? _GEN_2618 : _GEN_2986; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3052 = isAlloc_5 ? _GEN_2619 : _GEN_2987; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3053 = isAlloc_5 ? _GEN_2620 : _GEN_2988; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3054 = isAlloc_5 ? _GEN_2621 : _GEN_2989; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3055 = isAlloc_5 ? _GEN_2622 : _GEN_2990; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3056 = isAlloc_5 ? _GEN_2623 : _GEN_2991; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3057 = isAlloc_5 ? _GEN_2624 : _GEN_2992; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3058 = isAlloc_5 ? _GEN_2625 : _GEN_2993; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3059 = isAlloc_5 ? _GEN_2626 : _GEN_2994; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3060 = isAlloc_5 ? _GEN_2627 : _GEN_2995; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3061 = isAlloc_5 ? _GEN_2628 : _GEN_2996; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3062 = isAlloc_5 ? _GEN_2629 : _GEN_2997; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3063 = isAlloc_5 ? _GEN_2630 : _GEN_2998; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3064 = isAlloc_5 ? _GEN_2631 : _GEN_2999; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3065 = isAlloc_5 ? _GEN_2632 : _GEN_3000; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3066 = isAlloc_5 ? _GEN_2633 : _GEN_3001; // @[TBE.scala 109:24]
  wire  _GEN_3067 = isAlloc_5 ? _GEN_2634 : _GEN_2922; // @[TBE.scala 109:24]
  wire  _GEN_3068 = isAlloc_5 ? _GEN_2635 : _GEN_2923; // @[TBE.scala 109:24]
  wire  _GEN_3069 = isAlloc_5 ? _GEN_2636 : _GEN_2924; // @[TBE.scala 109:24]
  wire  _GEN_3070 = isAlloc_5 ? _GEN_2637 : _GEN_2925; // @[TBE.scala 109:24]
  wire  _GEN_3071 = isAlloc_5 ? _GEN_2638 : _GEN_2926; // @[TBE.scala 109:24]
  wire  _GEN_3072 = isAlloc_5 ? _GEN_2639 : _GEN_2927; // @[TBE.scala 109:24]
  wire  _GEN_3073 = isAlloc_5 ? _GEN_2640 : _GEN_2928; // @[TBE.scala 109:24]
  wire  _GEN_3074 = isAlloc_5 ? _GEN_2641 : _GEN_2929; // @[TBE.scala 109:24]
  wire  _GEN_3075 = isAlloc_5 ? _GEN_2642 : _GEN_2930; // @[TBE.scala 109:24]
  wire  _GEN_3076 = isAlloc_5 ? _GEN_2643 : _GEN_2931; // @[TBE.scala 109:24]
  wire  _GEN_3077 = isAlloc_5 ? _GEN_2644 : _GEN_2932; // @[TBE.scala 109:24]
  wire  _GEN_3078 = isAlloc_5 ? _GEN_2645 : _GEN_2933; // @[TBE.scala 109:24]
  wire  _GEN_3079 = isAlloc_5 ? _GEN_2646 : _GEN_2934; // @[TBE.scala 109:24]
  wire  _GEN_3080 = isAlloc_5 ? _GEN_2647 : _GEN_2935; // @[TBE.scala 109:24]
  wire  _GEN_3081 = isAlloc_5 ? _GEN_2648 : _GEN_2936; // @[TBE.scala 109:24]
  wire  _GEN_3082 = isAlloc_5 ? _GEN_2649 : _GEN_2937; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3084 = 4'h0 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3003; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3085 = 4'h1 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3004; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3086 = 4'h2 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3005; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3087 = 4'h3 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3006; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3088 = 4'h4 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3007; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3089 = 4'h5 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3008; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3090 = 4'h6 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3009; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3091 = 4'h7 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3010; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3092 = 4'h8 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3011; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3093 = 4'h9 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3012; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3094 = 4'ha == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3013; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3095 = 4'hb == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3014; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3096 = 4'hc == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3015; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3097 = 4'hd == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3016; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3098 = 4'he == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3017; // @[TBE.scala 110:27]
  wire [31:0] _GEN_3099 = 4'hf == idxAlloc[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3018; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3100 = 4'h0 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3019; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3101 = 4'h1 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3020; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3102 = 4'h2 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3021; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3103 = 4'h3 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3022; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3104 = 4'h4 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3023; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3105 = 4'h5 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3024; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3106 = 4'h6 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3025; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3107 = 4'h7 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3026; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3108 = 4'h8 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3027; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3109 = 4'h9 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3028; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3110 = 4'ha == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3029; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3111 = 4'hb == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3030; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3112 = 4'hc == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3031; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3113 = 4'hd == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3032; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3114 = 4'he == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3033; // @[TBE.scala 110:27]
  wire [2:0] _GEN_3115 = 4'hf == idxAlloc[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3034; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3116 = 4'h0 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3035; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3117 = 4'h1 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3036; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3118 = 4'h2 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3037; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3119 = 4'h3 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3038; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3120 = 4'h4 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3039; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3121 = 4'h5 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3040; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3122 = 4'h6 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3041; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3123 = 4'h7 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3042; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3124 = 4'h8 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3043; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3125 = 4'h9 == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3044; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3126 = 4'ha == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3045; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3127 = 4'hb == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3046; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3128 = 4'hc == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3047; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3129 = 4'hd == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3048; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3130 = 4'he == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3049; // @[TBE.scala 110:27]
  wire [1:0] _GEN_3131 = 4'hf == idxAlloc[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3050; // @[TBE.scala 110:27]
  wire  _GEN_3148 = _GEN_4161 | _GEN_3067; // @[TBE.scala 112:26]
  wire  _GEN_3149 = _GEN_4162 | _GEN_3068; // @[TBE.scala 112:26]
  wire  _GEN_3150 = _GEN_4163 | _GEN_3069; // @[TBE.scala 112:26]
  wire  _GEN_3151 = _GEN_4164 | _GEN_3070; // @[TBE.scala 112:26]
  wire  _GEN_3152 = _GEN_4165 | _GEN_3071; // @[TBE.scala 112:26]
  wire  _GEN_3153 = _GEN_4166 | _GEN_3072; // @[TBE.scala 112:26]
  wire  _GEN_3154 = _GEN_4167 | _GEN_3073; // @[TBE.scala 112:26]
  wire  _GEN_3155 = _GEN_4168 | _GEN_3074; // @[TBE.scala 112:26]
  wire  _GEN_3156 = _GEN_4169 | _GEN_3075; // @[TBE.scala 112:26]
  wire  _GEN_3157 = _GEN_4170 | _GEN_3076; // @[TBE.scala 112:26]
  wire  _GEN_3158 = _GEN_4171 | _GEN_3077; // @[TBE.scala 112:26]
  wire  _GEN_3159 = _GEN_4172 | _GEN_3078; // @[TBE.scala 112:26]
  wire  _GEN_3160 = _GEN_4173 | _GEN_3079; // @[TBE.scala 112:26]
  wire  _GEN_3161 = _GEN_4174 | _GEN_3080; // @[TBE.scala 112:26]
  wire  _GEN_3162 = _GEN_4175 | _GEN_3081; // @[TBE.scala 112:26]
  wire  _GEN_3163 = _GEN_4176 | _GEN_3082; // @[TBE.scala 112:26]
  wire  _T_301 = io_write_6_bits_command == 2'h2; // @[TBE.scala 137:46]
  wire  isDealloc_6 = _T_301 & io_write_6_valid; // @[TBE.scala 137:58]
  wire  _T_221 = isDealloc_6 & finder_6_io_value_valid; // @[TBE.scala 114:31]
  wire [4:0] idxUpdate_6 = {{1'd0}, finder_6_io_value_bits}; // @[TBE.scala 73:23 TBE.scala 104:18]
  wire  _GEN_3164 = 4'h0 == idxUpdate_6[3:0] ? 1'h0 : _GEN_3067; // @[TBE.scala 115:30]
  wire  _GEN_3165 = 4'h1 == idxUpdate_6[3:0] ? 1'h0 : _GEN_3068; // @[TBE.scala 115:30]
  wire  _GEN_3166 = 4'h2 == idxUpdate_6[3:0] ? 1'h0 : _GEN_3069; // @[TBE.scala 115:30]
  wire  _GEN_3167 = 4'h3 == idxUpdate_6[3:0] ? 1'h0 : _GEN_3070; // @[TBE.scala 115:30]
  wire  _GEN_3168 = 4'h4 == idxUpdate_6[3:0] ? 1'h0 : _GEN_3071; // @[TBE.scala 115:30]
  wire  _GEN_3169 = 4'h5 == idxUpdate_6[3:0] ? 1'h0 : _GEN_3072; // @[TBE.scala 115:30]
  wire  _GEN_3170 = 4'h6 == idxUpdate_6[3:0] ? 1'h0 : _GEN_3073; // @[TBE.scala 115:30]
  wire  _GEN_3171 = 4'h7 == idxUpdate_6[3:0] ? 1'h0 : _GEN_3074; // @[TBE.scala 115:30]
  wire  _GEN_3172 = 4'h8 == idxUpdate_6[3:0] ? 1'h0 : _GEN_3075; // @[TBE.scala 115:30]
  wire  _GEN_3173 = 4'h9 == idxUpdate_6[3:0] ? 1'h0 : _GEN_3076; // @[TBE.scala 115:30]
  wire  _GEN_3174 = 4'ha == idxUpdate_6[3:0] ? 1'h0 : _GEN_3077; // @[TBE.scala 115:30]
  wire  _GEN_3175 = 4'hb == idxUpdate_6[3:0] ? 1'h0 : _GEN_3078; // @[TBE.scala 115:30]
  wire  _GEN_3176 = 4'hc == idxUpdate_6[3:0] ? 1'h0 : _GEN_3079; // @[TBE.scala 115:30]
  wire  _GEN_3177 = 4'hd == idxUpdate_6[3:0] ? 1'h0 : _GEN_3080; // @[TBE.scala 115:30]
  wire  _GEN_3178 = 4'he == idxUpdate_6[3:0] ? 1'h0 : _GEN_3081; // @[TBE.scala 115:30]
  wire  _GEN_3179 = 4'hf == idxUpdate_6[3:0] ? 1'h0 : _GEN_3082; // @[TBE.scala 115:30]
  wire [31:0] _GEN_3180 = 4'h0 == idxUpdate_6[3:0] ? 32'h0 : _GEN_3003; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3181 = 4'h1 == idxUpdate_6[3:0] ? 32'h0 : _GEN_3004; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3182 = 4'h2 == idxUpdate_6[3:0] ? 32'h0 : _GEN_3005; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3183 = 4'h3 == idxUpdate_6[3:0] ? 32'h0 : _GEN_3006; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3184 = 4'h4 == idxUpdate_6[3:0] ? 32'h0 : _GEN_3007; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3185 = 4'h5 == idxUpdate_6[3:0] ? 32'h0 : _GEN_3008; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3186 = 4'h6 == idxUpdate_6[3:0] ? 32'h0 : _GEN_3009; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3187 = 4'h7 == idxUpdate_6[3:0] ? 32'h0 : _GEN_3010; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3188 = 4'h8 == idxUpdate_6[3:0] ? 32'h0 : _GEN_3011; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3189 = 4'h9 == idxUpdate_6[3:0] ? 32'h0 : _GEN_3012; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3190 = 4'ha == idxUpdate_6[3:0] ? 32'h0 : _GEN_3013; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3191 = 4'hb == idxUpdate_6[3:0] ? 32'h0 : _GEN_3014; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3192 = 4'hc == idxUpdate_6[3:0] ? 32'h0 : _GEN_3015; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3193 = 4'hd == idxUpdate_6[3:0] ? 32'h0 : _GEN_3016; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3194 = 4'he == idxUpdate_6[3:0] ? 32'h0 : _GEN_3017; // @[TBE.scala 116:31]
  wire [31:0] _GEN_3195 = 4'hf == idxUpdate_6[3:0] ? 32'h0 : _GEN_3018; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3196 = 4'h0 == idxUpdate_6[3:0] ? 3'h2 : _GEN_3019; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3197 = 4'h1 == idxUpdate_6[3:0] ? 3'h2 : _GEN_3020; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3198 = 4'h2 == idxUpdate_6[3:0] ? 3'h2 : _GEN_3021; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3199 = 4'h3 == idxUpdate_6[3:0] ? 3'h2 : _GEN_3022; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3200 = 4'h4 == idxUpdate_6[3:0] ? 3'h2 : _GEN_3023; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3201 = 4'h5 == idxUpdate_6[3:0] ? 3'h2 : _GEN_3024; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3202 = 4'h6 == idxUpdate_6[3:0] ? 3'h2 : _GEN_3025; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3203 = 4'h7 == idxUpdate_6[3:0] ? 3'h2 : _GEN_3026; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3204 = 4'h8 == idxUpdate_6[3:0] ? 3'h2 : _GEN_3027; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3205 = 4'h9 == idxUpdate_6[3:0] ? 3'h2 : _GEN_3028; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3206 = 4'ha == idxUpdate_6[3:0] ? 3'h2 : _GEN_3029; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3207 = 4'hb == idxUpdate_6[3:0] ? 3'h2 : _GEN_3030; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3208 = 4'hc == idxUpdate_6[3:0] ? 3'h2 : _GEN_3031; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3209 = 4'hd == idxUpdate_6[3:0] ? 3'h2 : _GEN_3032; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3210 = 4'he == idxUpdate_6[3:0] ? 3'h2 : _GEN_3033; // @[TBE.scala 116:31]
  wire [2:0] _GEN_3211 = 4'hf == idxUpdate_6[3:0] ? 3'h2 : _GEN_3034; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3212 = 4'h0 == idxUpdate_6[3:0] ? 2'h0 : _GEN_3035; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3213 = 4'h1 == idxUpdate_6[3:0] ? 2'h0 : _GEN_3036; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3214 = 4'h2 == idxUpdate_6[3:0] ? 2'h0 : _GEN_3037; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3215 = 4'h3 == idxUpdate_6[3:0] ? 2'h0 : _GEN_3038; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3216 = 4'h4 == idxUpdate_6[3:0] ? 2'h0 : _GEN_3039; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3217 = 4'h5 == idxUpdate_6[3:0] ? 2'h0 : _GEN_3040; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3218 = 4'h6 == idxUpdate_6[3:0] ? 2'h0 : _GEN_3041; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3219 = 4'h7 == idxUpdate_6[3:0] ? 2'h0 : _GEN_3042; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3220 = 4'h8 == idxUpdate_6[3:0] ? 2'h0 : _GEN_3043; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3221 = 4'h9 == idxUpdate_6[3:0] ? 2'h0 : _GEN_3044; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3222 = 4'ha == idxUpdate_6[3:0] ? 2'h0 : _GEN_3045; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3223 = 4'hb == idxUpdate_6[3:0] ? 2'h0 : _GEN_3046; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3224 = 4'hc == idxUpdate_6[3:0] ? 2'h0 : _GEN_3047; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3225 = 4'hd == idxUpdate_6[3:0] ? 2'h0 : _GEN_3048; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3226 = 4'he == idxUpdate_6[3:0] ? 2'h0 : _GEN_3049; // @[TBE.scala 116:31]
  wire [1:0] _GEN_3227 = 4'hf == idxUpdate_6[3:0] ? 2'h0 : _GEN_3050; // @[TBE.scala 116:31]
  wire  _T_303 = io_write_6_bits_command == 2'h3; // @[TBE.scala 138:44]
  wire  isWrite_6 = _T_303 & io_write_6_valid; // @[TBE.scala 138:55]
  wire  _T_229 = isWrite_6 & finder_6_io_value_valid; // @[TBE.scala 119:29]
  wire  _T_230 = ~io_write_6_bits_mask; // @[TBE.scala 120:35]
  wire [31:0] _GEN_3244 = 4'h0 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3003; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3245 = 4'h1 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3004; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3246 = 4'h2 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3005; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3247 = 4'h3 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3006; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3248 = 4'h4 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3007; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3249 = 4'h5 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3008; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3250 = 4'h6 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3009; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3251 = 4'h7 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3010; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3252 = 4'h8 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3011; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3253 = 4'h9 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3012; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3254 = 4'ha == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3013; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3255 = 4'hb == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3014; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3256 = 4'hc == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3015; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3257 = 4'hd == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3016; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3258 = 4'he == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3017; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3259 = 4'hf == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_fields_0 : _GEN_3018; // @[TBE.scala 121:63]
  wire [31:0] _GEN_3265 = 4'h1 == idxUpdate_6[3:0] ? TBEMemory_1_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3268 = 4'h2 == idxUpdate_6[3:0] ? TBEMemory_2_fields_0 : _GEN_3265; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3271 = 4'h3 == idxUpdate_6[3:0] ? TBEMemory_3_fields_0 : _GEN_3268; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3274 = 4'h4 == idxUpdate_6[3:0] ? TBEMemory_4_fields_0 : _GEN_3271; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3277 = 4'h5 == idxUpdate_6[3:0] ? TBEMemory_5_fields_0 : _GEN_3274; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3280 = 4'h6 == idxUpdate_6[3:0] ? TBEMemory_6_fields_0 : _GEN_3277; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3283 = 4'h7 == idxUpdate_6[3:0] ? TBEMemory_7_fields_0 : _GEN_3280; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3286 = 4'h8 == idxUpdate_6[3:0] ? TBEMemory_8_fields_0 : _GEN_3283; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3289 = 4'h9 == idxUpdate_6[3:0] ? TBEMemory_9_fields_0 : _GEN_3286; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3292 = 4'ha == idxUpdate_6[3:0] ? TBEMemory_10_fields_0 : _GEN_3289; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3295 = 4'hb == idxUpdate_6[3:0] ? TBEMemory_11_fields_0 : _GEN_3292; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3298 = 4'hc == idxUpdate_6[3:0] ? TBEMemory_12_fields_0 : _GEN_3295; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3301 = 4'hd == idxUpdate_6[3:0] ? TBEMemory_13_fields_0 : _GEN_3298; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3304 = 4'he == idxUpdate_6[3:0] ? TBEMemory_14_fields_0 : _GEN_3301; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3307 = 4'hf == idxUpdate_6[3:0] ? TBEMemory_15_fields_0 : _GEN_3304; // @[TBE.scala 122:15]
  wire [2:0] _GEN_3308 = 4'h0 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3019; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3309 = 4'h1 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3020; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3310 = 4'h2 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3021; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3311 = 4'h3 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3022; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3312 = 4'h4 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3023; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3313 = 4'h5 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3024; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3314 = 4'h6 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3025; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3315 = 4'h7 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3026; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3316 = 4'h8 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3027; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3317 = 4'h9 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3028; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3318 = 4'ha == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3029; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3319 = 4'hb == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3030; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3320 = 4'hc == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3031; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3321 = 4'hd == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3032; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3322 = 4'he == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3033; // @[TBE.scala 124:37]
  wire [2:0] _GEN_3323 = 4'hf == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_way : _GEN_3034; // @[TBE.scala 124:37]
  wire [1:0] _GEN_3324 = 4'h0 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3035; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3325 = 4'h1 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3036; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3326 = 4'h2 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3037; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3327 = 4'h3 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3038; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3328 = 4'h4 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3039; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3329 = 4'h5 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3040; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3330 = 4'h6 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3041; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3331 = 4'h7 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3042; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3332 = 4'h8 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3043; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3333 = 4'h9 == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3044; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3334 = 4'ha == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3045; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3335 = 4'hb == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3046; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3336 = 4'hc == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3047; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3337 = 4'hd == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3048; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3338 = 4'he == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3049; // @[TBE.scala 125:39]
  wire [1:0] _GEN_3339 = 4'hf == idxUpdate_6[3:0] ? io_write_6_bits_inputTBE_state_state : _GEN_3050; // @[TBE.scala 125:39]
  wire [31:0] _GEN_3340 = _T_230 ? _GEN_3244 : _GEN_3003; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3341 = _T_230 ? _GEN_3245 : _GEN_3004; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3342 = _T_230 ? _GEN_3246 : _GEN_3005; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3343 = _T_230 ? _GEN_3247 : _GEN_3006; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3344 = _T_230 ? _GEN_3248 : _GEN_3007; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3345 = _T_230 ? _GEN_3249 : _GEN_3008; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3346 = _T_230 ? _GEN_3250 : _GEN_3009; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3347 = _T_230 ? _GEN_3251 : _GEN_3010; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3348 = _T_230 ? _GEN_3252 : _GEN_3011; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3349 = _T_230 ? _GEN_3253 : _GEN_3012; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3350 = _T_230 ? _GEN_3254 : _GEN_3013; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3351 = _T_230 ? _GEN_3255 : _GEN_3014; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3352 = _T_230 ? _GEN_3256 : _GEN_3015; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3353 = _T_230 ? _GEN_3257 : _GEN_3016; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3354 = _T_230 ? _GEN_3258 : _GEN_3017; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3355 = _T_230 ? _GEN_3259 : _GEN_3018; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3356 = _T_230 ? _GEN_3019 : _GEN_3308; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3357 = _T_230 ? _GEN_3020 : _GEN_3309; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3358 = _T_230 ? _GEN_3021 : _GEN_3310; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3359 = _T_230 ? _GEN_3022 : _GEN_3311; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3360 = _T_230 ? _GEN_3023 : _GEN_3312; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3361 = _T_230 ? _GEN_3024 : _GEN_3313; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3362 = _T_230 ? _GEN_3025 : _GEN_3314; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3363 = _T_230 ? _GEN_3026 : _GEN_3315; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3364 = _T_230 ? _GEN_3027 : _GEN_3316; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3365 = _T_230 ? _GEN_3028 : _GEN_3317; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3366 = _T_230 ? _GEN_3029 : _GEN_3318; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3367 = _T_230 ? _GEN_3030 : _GEN_3319; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3368 = _T_230 ? _GEN_3031 : _GEN_3320; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3369 = _T_230 ? _GEN_3032 : _GEN_3321; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3370 = _T_230 ? _GEN_3033 : _GEN_3322; // @[TBE.scala 120:53]
  wire [2:0] _GEN_3371 = _T_230 ? _GEN_3034 : _GEN_3323; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3372 = _T_230 ? _GEN_3035 : _GEN_3324; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3373 = _T_230 ? _GEN_3036 : _GEN_3325; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3374 = _T_230 ? _GEN_3037 : _GEN_3326; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3375 = _T_230 ? _GEN_3038 : _GEN_3327; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3376 = _T_230 ? _GEN_3039 : _GEN_3328; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3377 = _T_230 ? _GEN_3040 : _GEN_3329; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3378 = _T_230 ? _GEN_3041 : _GEN_3330; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3379 = _T_230 ? _GEN_3042 : _GEN_3331; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3380 = _T_230 ? _GEN_3043 : _GEN_3332; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3381 = _T_230 ? _GEN_3044 : _GEN_3333; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3382 = _T_230 ? _GEN_3045 : _GEN_3334; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3383 = _T_230 ? _GEN_3046 : _GEN_3335; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3384 = _T_230 ? _GEN_3047 : _GEN_3336; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3385 = _T_230 ? _GEN_3048 : _GEN_3337; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3386 = _T_230 ? _GEN_3049 : _GEN_3338; // @[TBE.scala 120:53]
  wire [1:0] _GEN_3387 = _T_230 ? _GEN_3050 : _GEN_3339; // @[TBE.scala 120:53]
  wire [31:0] _GEN_3388 = _T_229 ? _GEN_3340 : _GEN_3003; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3389 = _T_229 ? _GEN_3341 : _GEN_3004; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3390 = _T_229 ? _GEN_3342 : _GEN_3005; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3391 = _T_229 ? _GEN_3343 : _GEN_3006; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3392 = _T_229 ? _GEN_3344 : _GEN_3007; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3393 = _T_229 ? _GEN_3345 : _GEN_3008; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3394 = _T_229 ? _GEN_3346 : _GEN_3009; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3395 = _T_229 ? _GEN_3347 : _GEN_3010; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3396 = _T_229 ? _GEN_3348 : _GEN_3011; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3397 = _T_229 ? _GEN_3349 : _GEN_3012; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3398 = _T_229 ? _GEN_3350 : _GEN_3013; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3399 = _T_229 ? _GEN_3351 : _GEN_3014; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3400 = _T_229 ? _GEN_3352 : _GEN_3015; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3401 = _T_229 ? _GEN_3353 : _GEN_3016; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3402 = _T_229 ? _GEN_3354 : _GEN_3017; // @[TBE.scala 119:57]
  wire [31:0] _GEN_3403 = _T_229 ? _GEN_3355 : _GEN_3018; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3404 = _T_229 ? _GEN_3356 : _GEN_3019; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3405 = _T_229 ? _GEN_3357 : _GEN_3020; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3406 = _T_229 ? _GEN_3358 : _GEN_3021; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3407 = _T_229 ? _GEN_3359 : _GEN_3022; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3408 = _T_229 ? _GEN_3360 : _GEN_3023; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3409 = _T_229 ? _GEN_3361 : _GEN_3024; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3410 = _T_229 ? _GEN_3362 : _GEN_3025; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3411 = _T_229 ? _GEN_3363 : _GEN_3026; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3412 = _T_229 ? _GEN_3364 : _GEN_3027; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3413 = _T_229 ? _GEN_3365 : _GEN_3028; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3414 = _T_229 ? _GEN_3366 : _GEN_3029; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3415 = _T_229 ? _GEN_3367 : _GEN_3030; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3416 = _T_229 ? _GEN_3368 : _GEN_3031; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3417 = _T_229 ? _GEN_3369 : _GEN_3032; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3418 = _T_229 ? _GEN_3370 : _GEN_3033; // @[TBE.scala 119:57]
  wire [2:0] _GEN_3419 = _T_229 ? _GEN_3371 : _GEN_3034; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3420 = _T_229 ? _GEN_3372 : _GEN_3035; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3421 = _T_229 ? _GEN_3373 : _GEN_3036; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3422 = _T_229 ? _GEN_3374 : _GEN_3037; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3423 = _T_229 ? _GEN_3375 : _GEN_3038; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3424 = _T_229 ? _GEN_3376 : _GEN_3039; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3425 = _T_229 ? _GEN_3377 : _GEN_3040; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3426 = _T_229 ? _GEN_3378 : _GEN_3041; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3427 = _T_229 ? _GEN_3379 : _GEN_3042; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3428 = _T_229 ? _GEN_3380 : _GEN_3043; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3429 = _T_229 ? _GEN_3381 : _GEN_3044; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3430 = _T_229 ? _GEN_3382 : _GEN_3045; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3431 = _T_229 ? _GEN_3383 : _GEN_3046; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3432 = _T_229 ? _GEN_3384 : _GEN_3047; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3433 = _T_229 ? _GEN_3385 : _GEN_3048; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3434 = _T_229 ? _GEN_3386 : _GEN_3049; // @[TBE.scala 119:57]
  wire [1:0] _GEN_3435 = _T_229 ? _GEN_3387 : _GEN_3050; // @[TBE.scala 119:57]
  wire  _GEN_3436 = _T_221 ? _GEN_3164 : _GEN_3067; // @[TBE.scala 114:59]
  wire  _GEN_3437 = _T_221 ? _GEN_3165 : _GEN_3068; // @[TBE.scala 114:59]
  wire  _GEN_3438 = _T_221 ? _GEN_3166 : _GEN_3069; // @[TBE.scala 114:59]
  wire  _GEN_3439 = _T_221 ? _GEN_3167 : _GEN_3070; // @[TBE.scala 114:59]
  wire  _GEN_3440 = _T_221 ? _GEN_3168 : _GEN_3071; // @[TBE.scala 114:59]
  wire  _GEN_3441 = _T_221 ? _GEN_3169 : _GEN_3072; // @[TBE.scala 114:59]
  wire  _GEN_3442 = _T_221 ? _GEN_3170 : _GEN_3073; // @[TBE.scala 114:59]
  wire  _GEN_3443 = _T_221 ? _GEN_3171 : _GEN_3074; // @[TBE.scala 114:59]
  wire  _GEN_3444 = _T_221 ? _GEN_3172 : _GEN_3075; // @[TBE.scala 114:59]
  wire  _GEN_3445 = _T_221 ? _GEN_3173 : _GEN_3076; // @[TBE.scala 114:59]
  wire  _GEN_3446 = _T_221 ? _GEN_3174 : _GEN_3077; // @[TBE.scala 114:59]
  wire  _GEN_3447 = _T_221 ? _GEN_3175 : _GEN_3078; // @[TBE.scala 114:59]
  wire  _GEN_3448 = _T_221 ? _GEN_3176 : _GEN_3079; // @[TBE.scala 114:59]
  wire  _GEN_3449 = _T_221 ? _GEN_3177 : _GEN_3080; // @[TBE.scala 114:59]
  wire  _GEN_3450 = _T_221 ? _GEN_3178 : _GEN_3081; // @[TBE.scala 114:59]
  wire  _GEN_3451 = _T_221 ? _GEN_3179 : _GEN_3082; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3452 = _T_221 ? _GEN_3180 : _GEN_3388; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3453 = _T_221 ? _GEN_3181 : _GEN_3389; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3454 = _T_221 ? _GEN_3182 : _GEN_3390; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3455 = _T_221 ? _GEN_3183 : _GEN_3391; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3456 = _T_221 ? _GEN_3184 : _GEN_3392; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3457 = _T_221 ? _GEN_3185 : _GEN_3393; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3458 = _T_221 ? _GEN_3186 : _GEN_3394; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3459 = _T_221 ? _GEN_3187 : _GEN_3395; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3460 = _T_221 ? _GEN_3188 : _GEN_3396; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3461 = _T_221 ? _GEN_3189 : _GEN_3397; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3462 = _T_221 ? _GEN_3190 : _GEN_3398; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3463 = _T_221 ? _GEN_3191 : _GEN_3399; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3464 = _T_221 ? _GEN_3192 : _GEN_3400; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3465 = _T_221 ? _GEN_3193 : _GEN_3401; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3466 = _T_221 ? _GEN_3194 : _GEN_3402; // @[TBE.scala 114:59]
  wire [31:0] _GEN_3467 = _T_221 ? _GEN_3195 : _GEN_3403; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3468 = _T_221 ? _GEN_3196 : _GEN_3404; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3469 = _T_221 ? _GEN_3197 : _GEN_3405; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3470 = _T_221 ? _GEN_3198 : _GEN_3406; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3471 = _T_221 ? _GEN_3199 : _GEN_3407; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3472 = _T_221 ? _GEN_3200 : _GEN_3408; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3473 = _T_221 ? _GEN_3201 : _GEN_3409; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3474 = _T_221 ? _GEN_3202 : _GEN_3410; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3475 = _T_221 ? _GEN_3203 : _GEN_3411; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3476 = _T_221 ? _GEN_3204 : _GEN_3412; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3477 = _T_221 ? _GEN_3205 : _GEN_3413; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3478 = _T_221 ? _GEN_3206 : _GEN_3414; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3479 = _T_221 ? _GEN_3207 : _GEN_3415; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3480 = _T_221 ? _GEN_3208 : _GEN_3416; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3481 = _T_221 ? _GEN_3209 : _GEN_3417; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3482 = _T_221 ? _GEN_3210 : _GEN_3418; // @[TBE.scala 114:59]
  wire [2:0] _GEN_3483 = _T_221 ? _GEN_3211 : _GEN_3419; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3484 = _T_221 ? _GEN_3212 : _GEN_3420; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3485 = _T_221 ? _GEN_3213 : _GEN_3421; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3486 = _T_221 ? _GEN_3214 : _GEN_3422; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3487 = _T_221 ? _GEN_3215 : _GEN_3423; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3488 = _T_221 ? _GEN_3216 : _GEN_3424; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3489 = _T_221 ? _GEN_3217 : _GEN_3425; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3490 = _T_221 ? _GEN_3218 : _GEN_3426; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3491 = _T_221 ? _GEN_3219 : _GEN_3427; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3492 = _T_221 ? _GEN_3220 : _GEN_3428; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3493 = _T_221 ? _GEN_3221 : _GEN_3429; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3494 = _T_221 ? _GEN_3222 : _GEN_3430; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3495 = _T_221 ? _GEN_3223 : _GEN_3431; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3496 = _T_221 ? _GEN_3224 : _GEN_3432; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3497 = _T_221 ? _GEN_3225 : _GEN_3433; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3498 = _T_221 ? _GEN_3226 : _GEN_3434; // @[TBE.scala 114:59]
  wire [1:0] _GEN_3499 = _T_221 ? _GEN_3227 : _GEN_3435; // @[TBE.scala 114:59]
  wire  _T_299 = io_write_6_bits_command == 2'h1; // @[TBE.scala 136:44]
  wire  isAlloc_6 = _T_299 & io_write_6_valid; // @[TBE.scala 136:54]
  wire [31:0] _GEN_3517 = isAlloc_6 ? _GEN_3084 : _GEN_3452; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3518 = isAlloc_6 ? _GEN_3085 : _GEN_3453; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3519 = isAlloc_6 ? _GEN_3086 : _GEN_3454; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3520 = isAlloc_6 ? _GEN_3087 : _GEN_3455; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3521 = isAlloc_6 ? _GEN_3088 : _GEN_3456; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3522 = isAlloc_6 ? _GEN_3089 : _GEN_3457; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3523 = isAlloc_6 ? _GEN_3090 : _GEN_3458; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3524 = isAlloc_6 ? _GEN_3091 : _GEN_3459; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3525 = isAlloc_6 ? _GEN_3092 : _GEN_3460; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3526 = isAlloc_6 ? _GEN_3093 : _GEN_3461; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3527 = isAlloc_6 ? _GEN_3094 : _GEN_3462; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3528 = isAlloc_6 ? _GEN_3095 : _GEN_3463; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3529 = isAlloc_6 ? _GEN_3096 : _GEN_3464; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3530 = isAlloc_6 ? _GEN_3097 : _GEN_3465; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3531 = isAlloc_6 ? _GEN_3098 : _GEN_3466; // @[TBE.scala 109:24]
  wire [31:0] _GEN_3532 = isAlloc_6 ? _GEN_3099 : _GEN_3467; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3533 = isAlloc_6 ? _GEN_3100 : _GEN_3468; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3534 = isAlloc_6 ? _GEN_3101 : _GEN_3469; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3535 = isAlloc_6 ? _GEN_3102 : _GEN_3470; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3536 = isAlloc_6 ? _GEN_3103 : _GEN_3471; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3537 = isAlloc_6 ? _GEN_3104 : _GEN_3472; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3538 = isAlloc_6 ? _GEN_3105 : _GEN_3473; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3539 = isAlloc_6 ? _GEN_3106 : _GEN_3474; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3540 = isAlloc_6 ? _GEN_3107 : _GEN_3475; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3541 = isAlloc_6 ? _GEN_3108 : _GEN_3476; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3542 = isAlloc_6 ? _GEN_3109 : _GEN_3477; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3543 = isAlloc_6 ? _GEN_3110 : _GEN_3478; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3544 = isAlloc_6 ? _GEN_3111 : _GEN_3479; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3545 = isAlloc_6 ? _GEN_3112 : _GEN_3480; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3546 = isAlloc_6 ? _GEN_3113 : _GEN_3481; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3547 = isAlloc_6 ? _GEN_3114 : _GEN_3482; // @[TBE.scala 109:24]
  wire [2:0] _GEN_3548 = isAlloc_6 ? _GEN_3115 : _GEN_3483; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3549 = isAlloc_6 ? _GEN_3116 : _GEN_3484; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3550 = isAlloc_6 ? _GEN_3117 : _GEN_3485; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3551 = isAlloc_6 ? _GEN_3118 : _GEN_3486; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3552 = isAlloc_6 ? _GEN_3119 : _GEN_3487; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3553 = isAlloc_6 ? _GEN_3120 : _GEN_3488; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3554 = isAlloc_6 ? _GEN_3121 : _GEN_3489; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3555 = isAlloc_6 ? _GEN_3122 : _GEN_3490; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3556 = isAlloc_6 ? _GEN_3123 : _GEN_3491; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3557 = isAlloc_6 ? _GEN_3124 : _GEN_3492; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3558 = isAlloc_6 ? _GEN_3125 : _GEN_3493; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3559 = isAlloc_6 ? _GEN_3126 : _GEN_3494; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3560 = isAlloc_6 ? _GEN_3127 : _GEN_3495; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3561 = isAlloc_6 ? _GEN_3128 : _GEN_3496; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3562 = isAlloc_6 ? _GEN_3129 : _GEN_3497; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3563 = isAlloc_6 ? _GEN_3130 : _GEN_3498; // @[TBE.scala 109:24]
  wire [1:0] _GEN_3564 = isAlloc_6 ? _GEN_3131 : _GEN_3499; // @[TBE.scala 109:24]
  wire  _GEN_3581 = isAlloc_6 ? _GEN_3148 : _GEN_3436; // @[TBE.scala 109:24]
  wire  _GEN_3582 = isAlloc_6 ? _GEN_3149 : _GEN_3437; // @[TBE.scala 109:24]
  wire  _GEN_3583 = isAlloc_6 ? _GEN_3150 : _GEN_3438; // @[TBE.scala 109:24]
  wire  _GEN_3584 = isAlloc_6 ? _GEN_3151 : _GEN_3439; // @[TBE.scala 109:24]
  wire  _GEN_3585 = isAlloc_6 ? _GEN_3152 : _GEN_3440; // @[TBE.scala 109:24]
  wire  _GEN_3586 = isAlloc_6 ? _GEN_3153 : _GEN_3441; // @[TBE.scala 109:24]
  wire  _GEN_3587 = isAlloc_6 ? _GEN_3154 : _GEN_3442; // @[TBE.scala 109:24]
  wire  _GEN_3588 = isAlloc_6 ? _GEN_3155 : _GEN_3443; // @[TBE.scala 109:24]
  wire  _GEN_3589 = isAlloc_6 ? _GEN_3156 : _GEN_3444; // @[TBE.scala 109:24]
  wire  _GEN_3590 = isAlloc_6 ? _GEN_3157 : _GEN_3445; // @[TBE.scala 109:24]
  wire  _GEN_3591 = isAlloc_6 ? _GEN_3158 : _GEN_3446; // @[TBE.scala 109:24]
  wire  _GEN_3592 = isAlloc_6 ? _GEN_3159 : _GEN_3447; // @[TBE.scala 109:24]
  wire  _GEN_3593 = isAlloc_6 ? _GEN_3160 : _GEN_3448; // @[TBE.scala 109:24]
  wire  _GEN_3594 = isAlloc_6 ? _GEN_3161 : _GEN_3449; // @[TBE.scala 109:24]
  wire  _GEN_3595 = isAlloc_6 ? _GEN_3162 : _GEN_3450; // @[TBE.scala 109:24]
  wire  _GEN_3596 = isAlloc_6 ? _GEN_3163 : _GEN_3451; // @[TBE.scala 109:24]
  wire  _GEN_3662 = _GEN_4161 | _GEN_3581; // @[TBE.scala 112:26]
  wire  _GEN_3663 = _GEN_4162 | _GEN_3582; // @[TBE.scala 112:26]
  wire  _GEN_3664 = _GEN_4163 | _GEN_3583; // @[TBE.scala 112:26]
  wire  _GEN_3665 = _GEN_4164 | _GEN_3584; // @[TBE.scala 112:26]
  wire  _GEN_3666 = _GEN_4165 | _GEN_3585; // @[TBE.scala 112:26]
  wire  _GEN_3667 = _GEN_4166 | _GEN_3586; // @[TBE.scala 112:26]
  wire  _GEN_3668 = _GEN_4167 | _GEN_3587; // @[TBE.scala 112:26]
  wire  _GEN_3669 = _GEN_4168 | _GEN_3588; // @[TBE.scala 112:26]
  wire  _GEN_3670 = _GEN_4169 | _GEN_3589; // @[TBE.scala 112:26]
  wire  _GEN_3671 = _GEN_4170 | _GEN_3590; // @[TBE.scala 112:26]
  wire  _GEN_3672 = _GEN_4171 | _GEN_3591; // @[TBE.scala 112:26]
  wire  _GEN_3673 = _GEN_4172 | _GEN_3592; // @[TBE.scala 112:26]
  wire  _GEN_3674 = _GEN_4173 | _GEN_3593; // @[TBE.scala 112:26]
  wire  _GEN_3675 = _GEN_4174 | _GEN_3594; // @[TBE.scala 112:26]
  wire  _GEN_3676 = _GEN_4175 | _GEN_3595; // @[TBE.scala 112:26]
  wire  _GEN_3677 = _GEN_4176 | _GEN_3596; // @[TBE.scala 112:26]
  wire  _T_307 = io_write_7_bits_command == 2'h2; // @[TBE.scala 137:46]
  wire  isDealloc_7 = _T_307 & io_write_7_valid; // @[TBE.scala 137:58]
  wire  _T_243 = isDealloc_7 & finder_7_io_value_valid; // @[TBE.scala 114:31]
  wire [4:0] idxUpdate_7 = {{1'd0}, finder_7_io_value_bits}; // @[TBE.scala 73:23 TBE.scala 104:18]
  wire  _T_309 = io_write_7_bits_command == 2'h3; // @[TBE.scala 138:44]
  wire  isWrite_7 = _T_309 & io_write_7_valid; // @[TBE.scala 138:55]
  wire  _T_251 = isWrite_7 & finder_7_io_value_valid; // @[TBE.scala 119:29]
  wire  _T_252 = ~io_write_7_bits_mask; // @[TBE.scala 120:35]
  wire [31:0] _GEN_3779 = 4'h1 == idxUpdate_7[3:0] ? TBEMemory_1_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3782 = 4'h2 == idxUpdate_7[3:0] ? TBEMemory_2_fields_0 : _GEN_3779; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3785 = 4'h3 == idxUpdate_7[3:0] ? TBEMemory_3_fields_0 : _GEN_3782; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3788 = 4'h4 == idxUpdate_7[3:0] ? TBEMemory_4_fields_0 : _GEN_3785; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3791 = 4'h5 == idxUpdate_7[3:0] ? TBEMemory_5_fields_0 : _GEN_3788; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3794 = 4'h6 == idxUpdate_7[3:0] ? TBEMemory_6_fields_0 : _GEN_3791; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3797 = 4'h7 == idxUpdate_7[3:0] ? TBEMemory_7_fields_0 : _GEN_3794; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3800 = 4'h8 == idxUpdate_7[3:0] ? TBEMemory_8_fields_0 : _GEN_3797; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3803 = 4'h9 == idxUpdate_7[3:0] ? TBEMemory_9_fields_0 : _GEN_3800; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3806 = 4'ha == idxUpdate_7[3:0] ? TBEMemory_10_fields_0 : _GEN_3803; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3809 = 4'hb == idxUpdate_7[3:0] ? TBEMemory_11_fields_0 : _GEN_3806; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3812 = 4'hc == idxUpdate_7[3:0] ? TBEMemory_12_fields_0 : _GEN_3809; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3815 = 4'hd == idxUpdate_7[3:0] ? TBEMemory_13_fields_0 : _GEN_3812; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3818 = 4'he == idxUpdate_7[3:0] ? TBEMemory_14_fields_0 : _GEN_3815; // @[TBE.scala 122:15]
  wire [31:0] _GEN_3821 = 4'hf == idxUpdate_7[3:0] ? TBEMemory_15_fields_0 : _GEN_3818; // @[TBE.scala 122:15]
  wire  _T_305 = io_write_7_bits_command == 2'h1; // @[TBE.scala 136:44]
  wire  isAlloc_7 = _T_305 & io_write_7_valid; // @[TBE.scala 136:54]
  wire [4:0] idxRead = {{1'd0}, finder_8_io_value_bits}; // @[TBE.scala 72:21 TBE.scala 95:11]
  wire [1:0] _GEN_4115 = 4'h1 == idxRead[3:0] ? TBEMemory_1_state_state : TBEMemory_0_state_state; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4116 = 4'h1 == idxRead[3:0] ? TBEMemory_1_way : TBEMemory_0_way; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4117 = 4'h1 == idxRead[3:0] ? TBEMemory_1_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4118 = 4'h2 == idxRead[3:0] ? TBEMemory_2_state_state : _GEN_4115; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4119 = 4'h2 == idxRead[3:0] ? TBEMemory_2_way : _GEN_4116; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4120 = 4'h2 == idxRead[3:0] ? TBEMemory_2_fields_0 : _GEN_4117; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4121 = 4'h3 == idxRead[3:0] ? TBEMemory_3_state_state : _GEN_4118; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4122 = 4'h3 == idxRead[3:0] ? TBEMemory_3_way : _GEN_4119; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4123 = 4'h3 == idxRead[3:0] ? TBEMemory_3_fields_0 : _GEN_4120; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4124 = 4'h4 == idxRead[3:0] ? TBEMemory_4_state_state : _GEN_4121; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4125 = 4'h4 == idxRead[3:0] ? TBEMemory_4_way : _GEN_4122; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4126 = 4'h4 == idxRead[3:0] ? TBEMemory_4_fields_0 : _GEN_4123; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4127 = 4'h5 == idxRead[3:0] ? TBEMemory_5_state_state : _GEN_4124; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4128 = 4'h5 == idxRead[3:0] ? TBEMemory_5_way : _GEN_4125; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4129 = 4'h5 == idxRead[3:0] ? TBEMemory_5_fields_0 : _GEN_4126; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4130 = 4'h6 == idxRead[3:0] ? TBEMemory_6_state_state : _GEN_4127; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4131 = 4'h6 == idxRead[3:0] ? TBEMemory_6_way : _GEN_4128; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4132 = 4'h6 == idxRead[3:0] ? TBEMemory_6_fields_0 : _GEN_4129; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4133 = 4'h7 == idxRead[3:0] ? TBEMemory_7_state_state : _GEN_4130; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4134 = 4'h7 == idxRead[3:0] ? TBEMemory_7_way : _GEN_4131; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4135 = 4'h7 == idxRead[3:0] ? TBEMemory_7_fields_0 : _GEN_4132; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4136 = 4'h8 == idxRead[3:0] ? TBEMemory_8_state_state : _GEN_4133; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4137 = 4'h8 == idxRead[3:0] ? TBEMemory_8_way : _GEN_4134; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4138 = 4'h8 == idxRead[3:0] ? TBEMemory_8_fields_0 : _GEN_4135; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4139 = 4'h9 == idxRead[3:0] ? TBEMemory_9_state_state : _GEN_4136; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4140 = 4'h9 == idxRead[3:0] ? TBEMemory_9_way : _GEN_4137; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4141 = 4'h9 == idxRead[3:0] ? TBEMemory_9_fields_0 : _GEN_4138; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4142 = 4'ha == idxRead[3:0] ? TBEMemory_10_state_state : _GEN_4139; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4143 = 4'ha == idxRead[3:0] ? TBEMemory_10_way : _GEN_4140; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4144 = 4'ha == idxRead[3:0] ? TBEMemory_10_fields_0 : _GEN_4141; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4145 = 4'hb == idxRead[3:0] ? TBEMemory_11_state_state : _GEN_4142; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4146 = 4'hb == idxRead[3:0] ? TBEMemory_11_way : _GEN_4143; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4147 = 4'hb == idxRead[3:0] ? TBEMemory_11_fields_0 : _GEN_4144; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4148 = 4'hc == idxRead[3:0] ? TBEMemory_12_state_state : _GEN_4145; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4149 = 4'hc == idxRead[3:0] ? TBEMemory_12_way : _GEN_4146; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4150 = 4'hc == idxRead[3:0] ? TBEMemory_12_fields_0 : _GEN_4147; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4151 = 4'hd == idxRead[3:0] ? TBEMemory_13_state_state : _GEN_4148; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4152 = 4'hd == idxRead[3:0] ? TBEMemory_13_way : _GEN_4149; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4153 = 4'hd == idxRead[3:0] ? TBEMemory_13_fields_0 : _GEN_4150; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4154 = 4'he == idxRead[3:0] ? TBEMemory_14_state_state : _GEN_4151; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4155 = 4'he == idxRead[3:0] ? TBEMemory_14_way : _GEN_4152; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4156 = 4'he == idxRead[3:0] ? TBEMemory_14_fields_0 : _GEN_4153; // @[TBE.scala 132:27]
  wire [1:0] _GEN_4157 = 4'hf == idxRead[3:0] ? TBEMemory_15_state_state : _GEN_4154; // @[TBE.scala 132:27]
  wire [2:0] _GEN_4158 = 4'hf == idxRead[3:0] ? TBEMemory_15_way : _GEN_4155; // @[TBE.scala 132:27]
  wire [31:0] _GEN_4159 = 4'hf == idxRead[3:0] ? TBEMemory_15_fields_0 : _GEN_4156; // @[TBE.scala 132:27]
  wire  _GEN_4289 = ~isAlloc_0; // @[TBE.scala 122:15]
  wire  _GEN_4290 = ~_T_89; // @[TBE.scala 122:15]
  wire  _GEN_4291 = _GEN_4289 & _GEN_4290; // @[TBE.scala 122:15]
  wire  _GEN_4292 = _GEN_4291 & _T_97; // @[TBE.scala 122:15]
  wire  _GEN_4293 = _GEN_4292 & _T_98; // @[TBE.scala 122:15]
  wire  _GEN_4294 = ~isAlloc_1; // @[TBE.scala 122:15]
  wire  _GEN_4295 = ~_T_111; // @[TBE.scala 122:15]
  wire  _GEN_4296 = _GEN_4294 & _GEN_4295; // @[TBE.scala 122:15]
  wire  _GEN_4297 = _GEN_4296 & _T_119; // @[TBE.scala 122:15]
  wire  _GEN_4298 = _GEN_4297 & _T_120; // @[TBE.scala 122:15]
  wire  _GEN_4299 = ~isAlloc_2; // @[TBE.scala 122:15]
  wire  _GEN_4300 = ~_T_133; // @[TBE.scala 122:15]
  wire  _GEN_4301 = _GEN_4299 & _GEN_4300; // @[TBE.scala 122:15]
  wire  _GEN_4302 = _GEN_4301 & _T_141; // @[TBE.scala 122:15]
  wire  _GEN_4303 = _GEN_4302 & _T_142; // @[TBE.scala 122:15]
  wire  _GEN_4304 = ~isAlloc_3; // @[TBE.scala 122:15]
  wire  _GEN_4305 = ~_T_155; // @[TBE.scala 122:15]
  wire  _GEN_4306 = _GEN_4304 & _GEN_4305; // @[TBE.scala 122:15]
  wire  _GEN_4307 = _GEN_4306 & _T_163; // @[TBE.scala 122:15]
  wire  _GEN_4308 = _GEN_4307 & _T_164; // @[TBE.scala 122:15]
  wire  _GEN_4309 = ~isAlloc_4; // @[TBE.scala 122:15]
  wire  _GEN_4310 = ~_T_177; // @[TBE.scala 122:15]
  wire  _GEN_4311 = _GEN_4309 & _GEN_4310; // @[TBE.scala 122:15]
  wire  _GEN_4312 = _GEN_4311 & _T_185; // @[TBE.scala 122:15]
  wire  _GEN_4313 = _GEN_4312 & _T_186; // @[TBE.scala 122:15]
  wire  _GEN_4314 = ~isAlloc_5; // @[TBE.scala 122:15]
  wire  _GEN_4315 = ~_T_199; // @[TBE.scala 122:15]
  wire  _GEN_4316 = _GEN_4314 & _GEN_4315; // @[TBE.scala 122:15]
  wire  _GEN_4317 = _GEN_4316 & _T_207; // @[TBE.scala 122:15]
  wire  _GEN_4318 = _GEN_4317 & _T_208; // @[TBE.scala 122:15]
  wire  _GEN_4319 = ~isAlloc_6; // @[TBE.scala 122:15]
  wire  _GEN_4320 = ~_T_221; // @[TBE.scala 122:15]
  wire  _GEN_4321 = _GEN_4319 & _GEN_4320; // @[TBE.scala 122:15]
  wire  _GEN_4322 = _GEN_4321 & _T_229; // @[TBE.scala 122:15]
  wire  _GEN_4323 = _GEN_4322 & _T_230; // @[TBE.scala 122:15]
  wire  _GEN_4324 = ~isAlloc_7; // @[TBE.scala 122:15]
  wire  _GEN_4325 = ~_T_243; // @[TBE.scala 122:15]
  wire  _GEN_4326 = _GEN_4324 & _GEN_4325; // @[TBE.scala 122:15]
  wire  _GEN_4327 = _GEN_4326 & _T_251; // @[TBE.scala 122:15]
  wire  _GEN_4328 = _GEN_4327 & _T_252; // @[TBE.scala 122:15]
  FindEmptyLine_9 allocLine ( // @[TBE.scala 79:25]
    .io_data_0(allocLine_io_data_0),
    .io_data_1(allocLine_io_data_1),
    .io_data_2(allocLine_io_data_2),
    .io_data_3(allocLine_io_data_3),
    .io_data_4(allocLine_io_data_4),
    .io_data_5(allocLine_io_data_5),
    .io_data_6(allocLine_io_data_6),
    .io_data_7(allocLine_io_data_7),
    .io_data_8(allocLine_io_data_8),
    .io_data_9(allocLine_io_data_9),
    .io_data_10(allocLine_io_data_10),
    .io_data_11(allocLine_io_data_11),
    .io_data_12(allocLine_io_data_12),
    .io_data_13(allocLine_io_data_13),
    .io_data_14(allocLine_io_data_14),
    .io_data_15(allocLine_io_data_15),
    .io_value_bits(allocLine_io_value_bits)
  );
  Find_9 finder_0 ( // @[TBE.scala 84:24]
    .io_key(finder_0_io_key),
    .io_data_0(finder_0_io_data_0),
    .io_data_1(finder_0_io_data_1),
    .io_data_2(finder_0_io_data_2),
    .io_data_3(finder_0_io_data_3),
    .io_data_4(finder_0_io_data_4),
    .io_data_5(finder_0_io_data_5),
    .io_data_6(finder_0_io_data_6),
    .io_data_7(finder_0_io_data_7),
    .io_data_8(finder_0_io_data_8),
    .io_data_9(finder_0_io_data_9),
    .io_data_10(finder_0_io_data_10),
    .io_data_11(finder_0_io_data_11),
    .io_data_12(finder_0_io_data_12),
    .io_data_13(finder_0_io_data_13),
    .io_data_14(finder_0_io_data_14),
    .io_data_15(finder_0_io_data_15),
    .io_valid_0(finder_0_io_valid_0),
    .io_valid_1(finder_0_io_valid_1),
    .io_valid_2(finder_0_io_valid_2),
    .io_valid_3(finder_0_io_valid_3),
    .io_valid_4(finder_0_io_valid_4),
    .io_valid_5(finder_0_io_valid_5),
    .io_valid_6(finder_0_io_valid_6),
    .io_valid_7(finder_0_io_valid_7),
    .io_valid_8(finder_0_io_valid_8),
    .io_valid_9(finder_0_io_valid_9),
    .io_valid_10(finder_0_io_valid_10),
    .io_valid_11(finder_0_io_valid_11),
    .io_valid_12(finder_0_io_valid_12),
    .io_valid_13(finder_0_io_valid_13),
    .io_valid_14(finder_0_io_valid_14),
    .io_valid_15(finder_0_io_valid_15),
    .io_value_valid(finder_0_io_value_valid),
    .io_value_bits(finder_0_io_value_bits)
  );
  Find_9 finder_1 ( // @[TBE.scala 84:24]
    .io_key(finder_1_io_key),
    .io_data_0(finder_1_io_data_0),
    .io_data_1(finder_1_io_data_1),
    .io_data_2(finder_1_io_data_2),
    .io_data_3(finder_1_io_data_3),
    .io_data_4(finder_1_io_data_4),
    .io_data_5(finder_1_io_data_5),
    .io_data_6(finder_1_io_data_6),
    .io_data_7(finder_1_io_data_7),
    .io_data_8(finder_1_io_data_8),
    .io_data_9(finder_1_io_data_9),
    .io_data_10(finder_1_io_data_10),
    .io_data_11(finder_1_io_data_11),
    .io_data_12(finder_1_io_data_12),
    .io_data_13(finder_1_io_data_13),
    .io_data_14(finder_1_io_data_14),
    .io_data_15(finder_1_io_data_15),
    .io_valid_0(finder_1_io_valid_0),
    .io_valid_1(finder_1_io_valid_1),
    .io_valid_2(finder_1_io_valid_2),
    .io_valid_3(finder_1_io_valid_3),
    .io_valid_4(finder_1_io_valid_4),
    .io_valid_5(finder_1_io_valid_5),
    .io_valid_6(finder_1_io_valid_6),
    .io_valid_7(finder_1_io_valid_7),
    .io_valid_8(finder_1_io_valid_8),
    .io_valid_9(finder_1_io_valid_9),
    .io_valid_10(finder_1_io_valid_10),
    .io_valid_11(finder_1_io_valid_11),
    .io_valid_12(finder_1_io_valid_12),
    .io_valid_13(finder_1_io_valid_13),
    .io_valid_14(finder_1_io_valid_14),
    .io_valid_15(finder_1_io_valid_15),
    .io_value_valid(finder_1_io_value_valid),
    .io_value_bits(finder_1_io_value_bits)
  );
  Find_9 finder_2 ( // @[TBE.scala 84:24]
    .io_key(finder_2_io_key),
    .io_data_0(finder_2_io_data_0),
    .io_data_1(finder_2_io_data_1),
    .io_data_2(finder_2_io_data_2),
    .io_data_3(finder_2_io_data_3),
    .io_data_4(finder_2_io_data_4),
    .io_data_5(finder_2_io_data_5),
    .io_data_6(finder_2_io_data_6),
    .io_data_7(finder_2_io_data_7),
    .io_data_8(finder_2_io_data_8),
    .io_data_9(finder_2_io_data_9),
    .io_data_10(finder_2_io_data_10),
    .io_data_11(finder_2_io_data_11),
    .io_data_12(finder_2_io_data_12),
    .io_data_13(finder_2_io_data_13),
    .io_data_14(finder_2_io_data_14),
    .io_data_15(finder_2_io_data_15),
    .io_valid_0(finder_2_io_valid_0),
    .io_valid_1(finder_2_io_valid_1),
    .io_valid_2(finder_2_io_valid_2),
    .io_valid_3(finder_2_io_valid_3),
    .io_valid_4(finder_2_io_valid_4),
    .io_valid_5(finder_2_io_valid_5),
    .io_valid_6(finder_2_io_valid_6),
    .io_valid_7(finder_2_io_valid_7),
    .io_valid_8(finder_2_io_valid_8),
    .io_valid_9(finder_2_io_valid_9),
    .io_valid_10(finder_2_io_valid_10),
    .io_valid_11(finder_2_io_valid_11),
    .io_valid_12(finder_2_io_valid_12),
    .io_valid_13(finder_2_io_valid_13),
    .io_valid_14(finder_2_io_valid_14),
    .io_valid_15(finder_2_io_valid_15),
    .io_value_valid(finder_2_io_value_valid),
    .io_value_bits(finder_2_io_value_bits)
  );
  Find_9 finder_3 ( // @[TBE.scala 84:24]
    .io_key(finder_3_io_key),
    .io_data_0(finder_3_io_data_0),
    .io_data_1(finder_3_io_data_1),
    .io_data_2(finder_3_io_data_2),
    .io_data_3(finder_3_io_data_3),
    .io_data_4(finder_3_io_data_4),
    .io_data_5(finder_3_io_data_5),
    .io_data_6(finder_3_io_data_6),
    .io_data_7(finder_3_io_data_7),
    .io_data_8(finder_3_io_data_8),
    .io_data_9(finder_3_io_data_9),
    .io_data_10(finder_3_io_data_10),
    .io_data_11(finder_3_io_data_11),
    .io_data_12(finder_3_io_data_12),
    .io_data_13(finder_3_io_data_13),
    .io_data_14(finder_3_io_data_14),
    .io_data_15(finder_3_io_data_15),
    .io_valid_0(finder_3_io_valid_0),
    .io_valid_1(finder_3_io_valid_1),
    .io_valid_2(finder_3_io_valid_2),
    .io_valid_3(finder_3_io_valid_3),
    .io_valid_4(finder_3_io_valid_4),
    .io_valid_5(finder_3_io_valid_5),
    .io_valid_6(finder_3_io_valid_6),
    .io_valid_7(finder_3_io_valid_7),
    .io_valid_8(finder_3_io_valid_8),
    .io_valid_9(finder_3_io_valid_9),
    .io_valid_10(finder_3_io_valid_10),
    .io_valid_11(finder_3_io_valid_11),
    .io_valid_12(finder_3_io_valid_12),
    .io_valid_13(finder_3_io_valid_13),
    .io_valid_14(finder_3_io_valid_14),
    .io_valid_15(finder_3_io_valid_15),
    .io_value_valid(finder_3_io_value_valid),
    .io_value_bits(finder_3_io_value_bits)
  );
  Find_9 finder_4 ( // @[TBE.scala 84:24]
    .io_key(finder_4_io_key),
    .io_data_0(finder_4_io_data_0),
    .io_data_1(finder_4_io_data_1),
    .io_data_2(finder_4_io_data_2),
    .io_data_3(finder_4_io_data_3),
    .io_data_4(finder_4_io_data_4),
    .io_data_5(finder_4_io_data_5),
    .io_data_6(finder_4_io_data_6),
    .io_data_7(finder_4_io_data_7),
    .io_data_8(finder_4_io_data_8),
    .io_data_9(finder_4_io_data_9),
    .io_data_10(finder_4_io_data_10),
    .io_data_11(finder_4_io_data_11),
    .io_data_12(finder_4_io_data_12),
    .io_data_13(finder_4_io_data_13),
    .io_data_14(finder_4_io_data_14),
    .io_data_15(finder_4_io_data_15),
    .io_valid_0(finder_4_io_valid_0),
    .io_valid_1(finder_4_io_valid_1),
    .io_valid_2(finder_4_io_valid_2),
    .io_valid_3(finder_4_io_valid_3),
    .io_valid_4(finder_4_io_valid_4),
    .io_valid_5(finder_4_io_valid_5),
    .io_valid_6(finder_4_io_valid_6),
    .io_valid_7(finder_4_io_valid_7),
    .io_valid_8(finder_4_io_valid_8),
    .io_valid_9(finder_4_io_valid_9),
    .io_valid_10(finder_4_io_valid_10),
    .io_valid_11(finder_4_io_valid_11),
    .io_valid_12(finder_4_io_valid_12),
    .io_valid_13(finder_4_io_valid_13),
    .io_valid_14(finder_4_io_valid_14),
    .io_valid_15(finder_4_io_valid_15),
    .io_value_valid(finder_4_io_value_valid),
    .io_value_bits(finder_4_io_value_bits)
  );
  Find_9 finder_5 ( // @[TBE.scala 84:24]
    .io_key(finder_5_io_key),
    .io_data_0(finder_5_io_data_0),
    .io_data_1(finder_5_io_data_1),
    .io_data_2(finder_5_io_data_2),
    .io_data_3(finder_5_io_data_3),
    .io_data_4(finder_5_io_data_4),
    .io_data_5(finder_5_io_data_5),
    .io_data_6(finder_5_io_data_6),
    .io_data_7(finder_5_io_data_7),
    .io_data_8(finder_5_io_data_8),
    .io_data_9(finder_5_io_data_9),
    .io_data_10(finder_5_io_data_10),
    .io_data_11(finder_5_io_data_11),
    .io_data_12(finder_5_io_data_12),
    .io_data_13(finder_5_io_data_13),
    .io_data_14(finder_5_io_data_14),
    .io_data_15(finder_5_io_data_15),
    .io_valid_0(finder_5_io_valid_0),
    .io_valid_1(finder_5_io_valid_1),
    .io_valid_2(finder_5_io_valid_2),
    .io_valid_3(finder_5_io_valid_3),
    .io_valid_4(finder_5_io_valid_4),
    .io_valid_5(finder_5_io_valid_5),
    .io_valid_6(finder_5_io_valid_6),
    .io_valid_7(finder_5_io_valid_7),
    .io_valid_8(finder_5_io_valid_8),
    .io_valid_9(finder_5_io_valid_9),
    .io_valid_10(finder_5_io_valid_10),
    .io_valid_11(finder_5_io_valid_11),
    .io_valid_12(finder_5_io_valid_12),
    .io_valid_13(finder_5_io_valid_13),
    .io_valid_14(finder_5_io_valid_14),
    .io_valid_15(finder_5_io_valid_15),
    .io_value_valid(finder_5_io_value_valid),
    .io_value_bits(finder_5_io_value_bits)
  );
  Find_9 finder_6 ( // @[TBE.scala 84:24]
    .io_key(finder_6_io_key),
    .io_data_0(finder_6_io_data_0),
    .io_data_1(finder_6_io_data_1),
    .io_data_2(finder_6_io_data_2),
    .io_data_3(finder_6_io_data_3),
    .io_data_4(finder_6_io_data_4),
    .io_data_5(finder_6_io_data_5),
    .io_data_6(finder_6_io_data_6),
    .io_data_7(finder_6_io_data_7),
    .io_data_8(finder_6_io_data_8),
    .io_data_9(finder_6_io_data_9),
    .io_data_10(finder_6_io_data_10),
    .io_data_11(finder_6_io_data_11),
    .io_data_12(finder_6_io_data_12),
    .io_data_13(finder_6_io_data_13),
    .io_data_14(finder_6_io_data_14),
    .io_data_15(finder_6_io_data_15),
    .io_valid_0(finder_6_io_valid_0),
    .io_valid_1(finder_6_io_valid_1),
    .io_valid_2(finder_6_io_valid_2),
    .io_valid_3(finder_6_io_valid_3),
    .io_valid_4(finder_6_io_valid_4),
    .io_valid_5(finder_6_io_valid_5),
    .io_valid_6(finder_6_io_valid_6),
    .io_valid_7(finder_6_io_valid_7),
    .io_valid_8(finder_6_io_valid_8),
    .io_valid_9(finder_6_io_valid_9),
    .io_valid_10(finder_6_io_valid_10),
    .io_valid_11(finder_6_io_valid_11),
    .io_valid_12(finder_6_io_valid_12),
    .io_valid_13(finder_6_io_valid_13),
    .io_valid_14(finder_6_io_valid_14),
    .io_valid_15(finder_6_io_valid_15),
    .io_value_valid(finder_6_io_value_valid),
    .io_value_bits(finder_6_io_value_bits)
  );
  Find_9 finder_7 ( // @[TBE.scala 84:24]
    .io_key(finder_7_io_key),
    .io_data_0(finder_7_io_data_0),
    .io_data_1(finder_7_io_data_1),
    .io_data_2(finder_7_io_data_2),
    .io_data_3(finder_7_io_data_3),
    .io_data_4(finder_7_io_data_4),
    .io_data_5(finder_7_io_data_5),
    .io_data_6(finder_7_io_data_6),
    .io_data_7(finder_7_io_data_7),
    .io_data_8(finder_7_io_data_8),
    .io_data_9(finder_7_io_data_9),
    .io_data_10(finder_7_io_data_10),
    .io_data_11(finder_7_io_data_11),
    .io_data_12(finder_7_io_data_12),
    .io_data_13(finder_7_io_data_13),
    .io_data_14(finder_7_io_data_14),
    .io_data_15(finder_7_io_data_15),
    .io_valid_0(finder_7_io_valid_0),
    .io_valid_1(finder_7_io_valid_1),
    .io_valid_2(finder_7_io_valid_2),
    .io_valid_3(finder_7_io_valid_3),
    .io_valid_4(finder_7_io_valid_4),
    .io_valid_5(finder_7_io_valid_5),
    .io_valid_6(finder_7_io_valid_6),
    .io_valid_7(finder_7_io_valid_7),
    .io_valid_8(finder_7_io_valid_8),
    .io_valid_9(finder_7_io_valid_9),
    .io_valid_10(finder_7_io_valid_10),
    .io_valid_11(finder_7_io_valid_11),
    .io_valid_12(finder_7_io_valid_12),
    .io_valid_13(finder_7_io_valid_13),
    .io_valid_14(finder_7_io_valid_14),
    .io_valid_15(finder_7_io_valid_15),
    .io_value_valid(finder_7_io_value_valid),
    .io_value_bits(finder_7_io_value_bits)
  );
  Find_9 finder_8 ( // @[TBE.scala 84:24]
    .io_key(finder_8_io_key),
    .io_data_0(finder_8_io_data_0),
    .io_data_1(finder_8_io_data_1),
    .io_data_2(finder_8_io_data_2),
    .io_data_3(finder_8_io_data_3),
    .io_data_4(finder_8_io_data_4),
    .io_data_5(finder_8_io_data_5),
    .io_data_6(finder_8_io_data_6),
    .io_data_7(finder_8_io_data_7),
    .io_data_8(finder_8_io_data_8),
    .io_data_9(finder_8_io_data_9),
    .io_data_10(finder_8_io_data_10),
    .io_data_11(finder_8_io_data_11),
    .io_data_12(finder_8_io_data_12),
    .io_data_13(finder_8_io_data_13),
    .io_data_14(finder_8_io_data_14),
    .io_data_15(finder_8_io_data_15),
    .io_valid_0(finder_8_io_valid_0),
    .io_valid_1(finder_8_io_valid_1),
    .io_valid_2(finder_8_io_valid_2),
    .io_valid_3(finder_8_io_valid_3),
    .io_valid_4(finder_8_io_valid_4),
    .io_valid_5(finder_8_io_valid_5),
    .io_valid_6(finder_8_io_valid_6),
    .io_valid_7(finder_8_io_valid_7),
    .io_valid_8(finder_8_io_valid_8),
    .io_valid_9(finder_8_io_valid_9),
    .io_valid_10(finder_8_io_valid_10),
    .io_valid_11(finder_8_io_valid_11),
    .io_valid_12(finder_8_io_valid_12),
    .io_valid_13(finder_8_io_valid_13),
    .io_valid_14(finder_8_io_valid_14),
    .io_valid_15(finder_8_io_valid_15),
    .io_value_valid(finder_8_io_value_valid),
    .io_value_bits(finder_8_io_value_bits)
  );
  assign io_outputTBE_bits_state_state = idxReadValid ? _GEN_4157 : 2'h0; // @[TBE.scala 132:21]
  assign io_outputTBE_bits_way = idxReadValid ? _GEN_4158 : 3'h2; // @[TBE.scala 132:21]
  assign io_outputTBE_bits_fields_0 = idxReadValid ? _GEN_4159 : 32'h0; // @[TBE.scala 132:21]
  assign io_isFull = _T_70 & _T_71; // @[TBE.scala 90:13]
  assign allocLine_io_data_0 = TBEValid_0; // @[TBE.scala 80:21]
  assign allocLine_io_data_1 = TBEValid_1; // @[TBE.scala 80:21]
  assign allocLine_io_data_2 = TBEValid_2; // @[TBE.scala 80:21]
  assign allocLine_io_data_3 = TBEValid_3; // @[TBE.scala 80:21]
  assign allocLine_io_data_4 = TBEValid_4; // @[TBE.scala 80:21]
  assign allocLine_io_data_5 = TBEValid_5; // @[TBE.scala 80:21]
  assign allocLine_io_data_6 = TBEValid_6; // @[TBE.scala 80:21]
  assign allocLine_io_data_7 = TBEValid_7; // @[TBE.scala 80:21]
  assign allocLine_io_data_8 = TBEValid_8; // @[TBE.scala 80:21]
  assign allocLine_io_data_9 = TBEValid_9; // @[TBE.scala 80:21]
  assign allocLine_io_data_10 = TBEValid_10; // @[TBE.scala 80:21]
  assign allocLine_io_data_11 = TBEValid_11; // @[TBE.scala 80:21]
  assign allocLine_io_data_12 = TBEValid_12; // @[TBE.scala 80:21]
  assign allocLine_io_data_13 = TBEValid_13; // @[TBE.scala 80:21]
  assign allocLine_io_data_14 = TBEValid_14; // @[TBE.scala 80:21]
  assign allocLine_io_data_15 = TBEValid_15; // @[TBE.scala 80:21]
  assign finder_0_io_key = io_write_0_bits_addr[31:0]; // @[TBE.scala 100:22]
  assign finder_0_io_data_0 = TBEAddr_0; // @[TBE.scala 101:23]
  assign finder_0_io_data_1 = TBEAddr_1; // @[TBE.scala 101:23]
  assign finder_0_io_data_2 = TBEAddr_2; // @[TBE.scala 101:23]
  assign finder_0_io_data_3 = TBEAddr_3; // @[TBE.scala 101:23]
  assign finder_0_io_data_4 = TBEAddr_4; // @[TBE.scala 101:23]
  assign finder_0_io_data_5 = TBEAddr_5; // @[TBE.scala 101:23]
  assign finder_0_io_data_6 = TBEAddr_6; // @[TBE.scala 101:23]
  assign finder_0_io_data_7 = TBEAddr_7; // @[TBE.scala 101:23]
  assign finder_0_io_data_8 = TBEAddr_8; // @[TBE.scala 101:23]
  assign finder_0_io_data_9 = TBEAddr_9; // @[TBE.scala 101:23]
  assign finder_0_io_data_10 = TBEAddr_10; // @[TBE.scala 101:23]
  assign finder_0_io_data_11 = TBEAddr_11; // @[TBE.scala 101:23]
  assign finder_0_io_data_12 = TBEAddr_12; // @[TBE.scala 101:23]
  assign finder_0_io_data_13 = TBEAddr_13; // @[TBE.scala 101:23]
  assign finder_0_io_data_14 = TBEAddr_14; // @[TBE.scala 101:23]
  assign finder_0_io_data_15 = TBEAddr_15; // @[TBE.scala 101:23]
  assign finder_0_io_valid_0 = TBEValid_0; // @[TBE.scala 102:24]
  assign finder_0_io_valid_1 = TBEValid_1; // @[TBE.scala 102:24]
  assign finder_0_io_valid_2 = TBEValid_2; // @[TBE.scala 102:24]
  assign finder_0_io_valid_3 = TBEValid_3; // @[TBE.scala 102:24]
  assign finder_0_io_valid_4 = TBEValid_4; // @[TBE.scala 102:24]
  assign finder_0_io_valid_5 = TBEValid_5; // @[TBE.scala 102:24]
  assign finder_0_io_valid_6 = TBEValid_6; // @[TBE.scala 102:24]
  assign finder_0_io_valid_7 = TBEValid_7; // @[TBE.scala 102:24]
  assign finder_0_io_valid_8 = TBEValid_8; // @[TBE.scala 102:24]
  assign finder_0_io_valid_9 = TBEValid_9; // @[TBE.scala 102:24]
  assign finder_0_io_valid_10 = TBEValid_10; // @[TBE.scala 102:24]
  assign finder_0_io_valid_11 = TBEValid_11; // @[TBE.scala 102:24]
  assign finder_0_io_valid_12 = TBEValid_12; // @[TBE.scala 102:24]
  assign finder_0_io_valid_13 = TBEValid_13; // @[TBE.scala 102:24]
  assign finder_0_io_valid_14 = TBEValid_14; // @[TBE.scala 102:24]
  assign finder_0_io_valid_15 = TBEValid_15; // @[TBE.scala 102:24]
  assign finder_1_io_key = io_write_1_bits_addr[31:0]; // @[TBE.scala 100:22]
  assign finder_1_io_data_0 = TBEAddr_0; // @[TBE.scala 101:23]
  assign finder_1_io_data_1 = TBEAddr_1; // @[TBE.scala 101:23]
  assign finder_1_io_data_2 = TBEAddr_2; // @[TBE.scala 101:23]
  assign finder_1_io_data_3 = TBEAddr_3; // @[TBE.scala 101:23]
  assign finder_1_io_data_4 = TBEAddr_4; // @[TBE.scala 101:23]
  assign finder_1_io_data_5 = TBEAddr_5; // @[TBE.scala 101:23]
  assign finder_1_io_data_6 = TBEAddr_6; // @[TBE.scala 101:23]
  assign finder_1_io_data_7 = TBEAddr_7; // @[TBE.scala 101:23]
  assign finder_1_io_data_8 = TBEAddr_8; // @[TBE.scala 101:23]
  assign finder_1_io_data_9 = TBEAddr_9; // @[TBE.scala 101:23]
  assign finder_1_io_data_10 = TBEAddr_10; // @[TBE.scala 101:23]
  assign finder_1_io_data_11 = TBEAddr_11; // @[TBE.scala 101:23]
  assign finder_1_io_data_12 = TBEAddr_12; // @[TBE.scala 101:23]
  assign finder_1_io_data_13 = TBEAddr_13; // @[TBE.scala 101:23]
  assign finder_1_io_data_14 = TBEAddr_14; // @[TBE.scala 101:23]
  assign finder_1_io_data_15 = TBEAddr_15; // @[TBE.scala 101:23]
  assign finder_1_io_valid_0 = TBEValid_0; // @[TBE.scala 102:24]
  assign finder_1_io_valid_1 = TBEValid_1; // @[TBE.scala 102:24]
  assign finder_1_io_valid_2 = TBEValid_2; // @[TBE.scala 102:24]
  assign finder_1_io_valid_3 = TBEValid_3; // @[TBE.scala 102:24]
  assign finder_1_io_valid_4 = TBEValid_4; // @[TBE.scala 102:24]
  assign finder_1_io_valid_5 = TBEValid_5; // @[TBE.scala 102:24]
  assign finder_1_io_valid_6 = TBEValid_6; // @[TBE.scala 102:24]
  assign finder_1_io_valid_7 = TBEValid_7; // @[TBE.scala 102:24]
  assign finder_1_io_valid_8 = TBEValid_8; // @[TBE.scala 102:24]
  assign finder_1_io_valid_9 = TBEValid_9; // @[TBE.scala 102:24]
  assign finder_1_io_valid_10 = TBEValid_10; // @[TBE.scala 102:24]
  assign finder_1_io_valid_11 = TBEValid_11; // @[TBE.scala 102:24]
  assign finder_1_io_valid_12 = TBEValid_12; // @[TBE.scala 102:24]
  assign finder_1_io_valid_13 = TBEValid_13; // @[TBE.scala 102:24]
  assign finder_1_io_valid_14 = TBEValid_14; // @[TBE.scala 102:24]
  assign finder_1_io_valid_15 = TBEValid_15; // @[TBE.scala 102:24]
  assign finder_2_io_key = io_write_2_bits_addr[31:0]; // @[TBE.scala 100:22]
  assign finder_2_io_data_0 = TBEAddr_0; // @[TBE.scala 101:23]
  assign finder_2_io_data_1 = TBEAddr_1; // @[TBE.scala 101:23]
  assign finder_2_io_data_2 = TBEAddr_2; // @[TBE.scala 101:23]
  assign finder_2_io_data_3 = TBEAddr_3; // @[TBE.scala 101:23]
  assign finder_2_io_data_4 = TBEAddr_4; // @[TBE.scala 101:23]
  assign finder_2_io_data_5 = TBEAddr_5; // @[TBE.scala 101:23]
  assign finder_2_io_data_6 = TBEAddr_6; // @[TBE.scala 101:23]
  assign finder_2_io_data_7 = TBEAddr_7; // @[TBE.scala 101:23]
  assign finder_2_io_data_8 = TBEAddr_8; // @[TBE.scala 101:23]
  assign finder_2_io_data_9 = TBEAddr_9; // @[TBE.scala 101:23]
  assign finder_2_io_data_10 = TBEAddr_10; // @[TBE.scala 101:23]
  assign finder_2_io_data_11 = TBEAddr_11; // @[TBE.scala 101:23]
  assign finder_2_io_data_12 = TBEAddr_12; // @[TBE.scala 101:23]
  assign finder_2_io_data_13 = TBEAddr_13; // @[TBE.scala 101:23]
  assign finder_2_io_data_14 = TBEAddr_14; // @[TBE.scala 101:23]
  assign finder_2_io_data_15 = TBEAddr_15; // @[TBE.scala 101:23]
  assign finder_2_io_valid_0 = TBEValid_0; // @[TBE.scala 102:24]
  assign finder_2_io_valid_1 = TBEValid_1; // @[TBE.scala 102:24]
  assign finder_2_io_valid_2 = TBEValid_2; // @[TBE.scala 102:24]
  assign finder_2_io_valid_3 = TBEValid_3; // @[TBE.scala 102:24]
  assign finder_2_io_valid_4 = TBEValid_4; // @[TBE.scala 102:24]
  assign finder_2_io_valid_5 = TBEValid_5; // @[TBE.scala 102:24]
  assign finder_2_io_valid_6 = TBEValid_6; // @[TBE.scala 102:24]
  assign finder_2_io_valid_7 = TBEValid_7; // @[TBE.scala 102:24]
  assign finder_2_io_valid_8 = TBEValid_8; // @[TBE.scala 102:24]
  assign finder_2_io_valid_9 = TBEValid_9; // @[TBE.scala 102:24]
  assign finder_2_io_valid_10 = TBEValid_10; // @[TBE.scala 102:24]
  assign finder_2_io_valid_11 = TBEValid_11; // @[TBE.scala 102:24]
  assign finder_2_io_valid_12 = TBEValid_12; // @[TBE.scala 102:24]
  assign finder_2_io_valid_13 = TBEValid_13; // @[TBE.scala 102:24]
  assign finder_2_io_valid_14 = TBEValid_14; // @[TBE.scala 102:24]
  assign finder_2_io_valid_15 = TBEValid_15; // @[TBE.scala 102:24]
  assign finder_3_io_key = io_write_3_bits_addr[31:0]; // @[TBE.scala 100:22]
  assign finder_3_io_data_0 = TBEAddr_0; // @[TBE.scala 101:23]
  assign finder_3_io_data_1 = TBEAddr_1; // @[TBE.scala 101:23]
  assign finder_3_io_data_2 = TBEAddr_2; // @[TBE.scala 101:23]
  assign finder_3_io_data_3 = TBEAddr_3; // @[TBE.scala 101:23]
  assign finder_3_io_data_4 = TBEAddr_4; // @[TBE.scala 101:23]
  assign finder_3_io_data_5 = TBEAddr_5; // @[TBE.scala 101:23]
  assign finder_3_io_data_6 = TBEAddr_6; // @[TBE.scala 101:23]
  assign finder_3_io_data_7 = TBEAddr_7; // @[TBE.scala 101:23]
  assign finder_3_io_data_8 = TBEAddr_8; // @[TBE.scala 101:23]
  assign finder_3_io_data_9 = TBEAddr_9; // @[TBE.scala 101:23]
  assign finder_3_io_data_10 = TBEAddr_10; // @[TBE.scala 101:23]
  assign finder_3_io_data_11 = TBEAddr_11; // @[TBE.scala 101:23]
  assign finder_3_io_data_12 = TBEAddr_12; // @[TBE.scala 101:23]
  assign finder_3_io_data_13 = TBEAddr_13; // @[TBE.scala 101:23]
  assign finder_3_io_data_14 = TBEAddr_14; // @[TBE.scala 101:23]
  assign finder_3_io_data_15 = TBEAddr_15; // @[TBE.scala 101:23]
  assign finder_3_io_valid_0 = TBEValid_0; // @[TBE.scala 102:24]
  assign finder_3_io_valid_1 = TBEValid_1; // @[TBE.scala 102:24]
  assign finder_3_io_valid_2 = TBEValid_2; // @[TBE.scala 102:24]
  assign finder_3_io_valid_3 = TBEValid_3; // @[TBE.scala 102:24]
  assign finder_3_io_valid_4 = TBEValid_4; // @[TBE.scala 102:24]
  assign finder_3_io_valid_5 = TBEValid_5; // @[TBE.scala 102:24]
  assign finder_3_io_valid_6 = TBEValid_6; // @[TBE.scala 102:24]
  assign finder_3_io_valid_7 = TBEValid_7; // @[TBE.scala 102:24]
  assign finder_3_io_valid_8 = TBEValid_8; // @[TBE.scala 102:24]
  assign finder_3_io_valid_9 = TBEValid_9; // @[TBE.scala 102:24]
  assign finder_3_io_valid_10 = TBEValid_10; // @[TBE.scala 102:24]
  assign finder_3_io_valid_11 = TBEValid_11; // @[TBE.scala 102:24]
  assign finder_3_io_valid_12 = TBEValid_12; // @[TBE.scala 102:24]
  assign finder_3_io_valid_13 = TBEValid_13; // @[TBE.scala 102:24]
  assign finder_3_io_valid_14 = TBEValid_14; // @[TBE.scala 102:24]
  assign finder_3_io_valid_15 = TBEValid_15; // @[TBE.scala 102:24]
  assign finder_4_io_key = io_write_4_bits_addr[31:0]; // @[TBE.scala 100:22]
  assign finder_4_io_data_0 = TBEAddr_0; // @[TBE.scala 101:23]
  assign finder_4_io_data_1 = TBEAddr_1; // @[TBE.scala 101:23]
  assign finder_4_io_data_2 = TBEAddr_2; // @[TBE.scala 101:23]
  assign finder_4_io_data_3 = TBEAddr_3; // @[TBE.scala 101:23]
  assign finder_4_io_data_4 = TBEAddr_4; // @[TBE.scala 101:23]
  assign finder_4_io_data_5 = TBEAddr_5; // @[TBE.scala 101:23]
  assign finder_4_io_data_6 = TBEAddr_6; // @[TBE.scala 101:23]
  assign finder_4_io_data_7 = TBEAddr_7; // @[TBE.scala 101:23]
  assign finder_4_io_data_8 = TBEAddr_8; // @[TBE.scala 101:23]
  assign finder_4_io_data_9 = TBEAddr_9; // @[TBE.scala 101:23]
  assign finder_4_io_data_10 = TBEAddr_10; // @[TBE.scala 101:23]
  assign finder_4_io_data_11 = TBEAddr_11; // @[TBE.scala 101:23]
  assign finder_4_io_data_12 = TBEAddr_12; // @[TBE.scala 101:23]
  assign finder_4_io_data_13 = TBEAddr_13; // @[TBE.scala 101:23]
  assign finder_4_io_data_14 = TBEAddr_14; // @[TBE.scala 101:23]
  assign finder_4_io_data_15 = TBEAddr_15; // @[TBE.scala 101:23]
  assign finder_4_io_valid_0 = TBEValid_0; // @[TBE.scala 102:24]
  assign finder_4_io_valid_1 = TBEValid_1; // @[TBE.scala 102:24]
  assign finder_4_io_valid_2 = TBEValid_2; // @[TBE.scala 102:24]
  assign finder_4_io_valid_3 = TBEValid_3; // @[TBE.scala 102:24]
  assign finder_4_io_valid_4 = TBEValid_4; // @[TBE.scala 102:24]
  assign finder_4_io_valid_5 = TBEValid_5; // @[TBE.scala 102:24]
  assign finder_4_io_valid_6 = TBEValid_6; // @[TBE.scala 102:24]
  assign finder_4_io_valid_7 = TBEValid_7; // @[TBE.scala 102:24]
  assign finder_4_io_valid_8 = TBEValid_8; // @[TBE.scala 102:24]
  assign finder_4_io_valid_9 = TBEValid_9; // @[TBE.scala 102:24]
  assign finder_4_io_valid_10 = TBEValid_10; // @[TBE.scala 102:24]
  assign finder_4_io_valid_11 = TBEValid_11; // @[TBE.scala 102:24]
  assign finder_4_io_valid_12 = TBEValid_12; // @[TBE.scala 102:24]
  assign finder_4_io_valid_13 = TBEValid_13; // @[TBE.scala 102:24]
  assign finder_4_io_valid_14 = TBEValid_14; // @[TBE.scala 102:24]
  assign finder_4_io_valid_15 = TBEValid_15; // @[TBE.scala 102:24]
  assign finder_5_io_key = io_write_5_bits_addr[31:0]; // @[TBE.scala 100:22]
  assign finder_5_io_data_0 = TBEAddr_0; // @[TBE.scala 101:23]
  assign finder_5_io_data_1 = TBEAddr_1; // @[TBE.scala 101:23]
  assign finder_5_io_data_2 = TBEAddr_2; // @[TBE.scala 101:23]
  assign finder_5_io_data_3 = TBEAddr_3; // @[TBE.scala 101:23]
  assign finder_5_io_data_4 = TBEAddr_4; // @[TBE.scala 101:23]
  assign finder_5_io_data_5 = TBEAddr_5; // @[TBE.scala 101:23]
  assign finder_5_io_data_6 = TBEAddr_6; // @[TBE.scala 101:23]
  assign finder_5_io_data_7 = TBEAddr_7; // @[TBE.scala 101:23]
  assign finder_5_io_data_8 = TBEAddr_8; // @[TBE.scala 101:23]
  assign finder_5_io_data_9 = TBEAddr_9; // @[TBE.scala 101:23]
  assign finder_5_io_data_10 = TBEAddr_10; // @[TBE.scala 101:23]
  assign finder_5_io_data_11 = TBEAddr_11; // @[TBE.scala 101:23]
  assign finder_5_io_data_12 = TBEAddr_12; // @[TBE.scala 101:23]
  assign finder_5_io_data_13 = TBEAddr_13; // @[TBE.scala 101:23]
  assign finder_5_io_data_14 = TBEAddr_14; // @[TBE.scala 101:23]
  assign finder_5_io_data_15 = TBEAddr_15; // @[TBE.scala 101:23]
  assign finder_5_io_valid_0 = TBEValid_0; // @[TBE.scala 102:24]
  assign finder_5_io_valid_1 = TBEValid_1; // @[TBE.scala 102:24]
  assign finder_5_io_valid_2 = TBEValid_2; // @[TBE.scala 102:24]
  assign finder_5_io_valid_3 = TBEValid_3; // @[TBE.scala 102:24]
  assign finder_5_io_valid_4 = TBEValid_4; // @[TBE.scala 102:24]
  assign finder_5_io_valid_5 = TBEValid_5; // @[TBE.scala 102:24]
  assign finder_5_io_valid_6 = TBEValid_6; // @[TBE.scala 102:24]
  assign finder_5_io_valid_7 = TBEValid_7; // @[TBE.scala 102:24]
  assign finder_5_io_valid_8 = TBEValid_8; // @[TBE.scala 102:24]
  assign finder_5_io_valid_9 = TBEValid_9; // @[TBE.scala 102:24]
  assign finder_5_io_valid_10 = TBEValid_10; // @[TBE.scala 102:24]
  assign finder_5_io_valid_11 = TBEValid_11; // @[TBE.scala 102:24]
  assign finder_5_io_valid_12 = TBEValid_12; // @[TBE.scala 102:24]
  assign finder_5_io_valid_13 = TBEValid_13; // @[TBE.scala 102:24]
  assign finder_5_io_valid_14 = TBEValid_14; // @[TBE.scala 102:24]
  assign finder_5_io_valid_15 = TBEValid_15; // @[TBE.scala 102:24]
  assign finder_6_io_key = io_write_6_bits_addr[31:0]; // @[TBE.scala 100:22]
  assign finder_6_io_data_0 = TBEAddr_0; // @[TBE.scala 101:23]
  assign finder_6_io_data_1 = TBEAddr_1; // @[TBE.scala 101:23]
  assign finder_6_io_data_2 = TBEAddr_2; // @[TBE.scala 101:23]
  assign finder_6_io_data_3 = TBEAddr_3; // @[TBE.scala 101:23]
  assign finder_6_io_data_4 = TBEAddr_4; // @[TBE.scala 101:23]
  assign finder_6_io_data_5 = TBEAddr_5; // @[TBE.scala 101:23]
  assign finder_6_io_data_6 = TBEAddr_6; // @[TBE.scala 101:23]
  assign finder_6_io_data_7 = TBEAddr_7; // @[TBE.scala 101:23]
  assign finder_6_io_data_8 = TBEAddr_8; // @[TBE.scala 101:23]
  assign finder_6_io_data_9 = TBEAddr_9; // @[TBE.scala 101:23]
  assign finder_6_io_data_10 = TBEAddr_10; // @[TBE.scala 101:23]
  assign finder_6_io_data_11 = TBEAddr_11; // @[TBE.scala 101:23]
  assign finder_6_io_data_12 = TBEAddr_12; // @[TBE.scala 101:23]
  assign finder_6_io_data_13 = TBEAddr_13; // @[TBE.scala 101:23]
  assign finder_6_io_data_14 = TBEAddr_14; // @[TBE.scala 101:23]
  assign finder_6_io_data_15 = TBEAddr_15; // @[TBE.scala 101:23]
  assign finder_6_io_valid_0 = TBEValid_0; // @[TBE.scala 102:24]
  assign finder_6_io_valid_1 = TBEValid_1; // @[TBE.scala 102:24]
  assign finder_6_io_valid_2 = TBEValid_2; // @[TBE.scala 102:24]
  assign finder_6_io_valid_3 = TBEValid_3; // @[TBE.scala 102:24]
  assign finder_6_io_valid_4 = TBEValid_4; // @[TBE.scala 102:24]
  assign finder_6_io_valid_5 = TBEValid_5; // @[TBE.scala 102:24]
  assign finder_6_io_valid_6 = TBEValid_6; // @[TBE.scala 102:24]
  assign finder_6_io_valid_7 = TBEValid_7; // @[TBE.scala 102:24]
  assign finder_6_io_valid_8 = TBEValid_8; // @[TBE.scala 102:24]
  assign finder_6_io_valid_9 = TBEValid_9; // @[TBE.scala 102:24]
  assign finder_6_io_valid_10 = TBEValid_10; // @[TBE.scala 102:24]
  assign finder_6_io_valid_11 = TBEValid_11; // @[TBE.scala 102:24]
  assign finder_6_io_valid_12 = TBEValid_12; // @[TBE.scala 102:24]
  assign finder_6_io_valid_13 = TBEValid_13; // @[TBE.scala 102:24]
  assign finder_6_io_valid_14 = TBEValid_14; // @[TBE.scala 102:24]
  assign finder_6_io_valid_15 = TBEValid_15; // @[TBE.scala 102:24]
  assign finder_7_io_key = io_write_7_bits_addr[31:0]; // @[TBE.scala 100:22]
  assign finder_7_io_data_0 = TBEAddr_0; // @[TBE.scala 101:23]
  assign finder_7_io_data_1 = TBEAddr_1; // @[TBE.scala 101:23]
  assign finder_7_io_data_2 = TBEAddr_2; // @[TBE.scala 101:23]
  assign finder_7_io_data_3 = TBEAddr_3; // @[TBE.scala 101:23]
  assign finder_7_io_data_4 = TBEAddr_4; // @[TBE.scala 101:23]
  assign finder_7_io_data_5 = TBEAddr_5; // @[TBE.scala 101:23]
  assign finder_7_io_data_6 = TBEAddr_6; // @[TBE.scala 101:23]
  assign finder_7_io_data_7 = TBEAddr_7; // @[TBE.scala 101:23]
  assign finder_7_io_data_8 = TBEAddr_8; // @[TBE.scala 101:23]
  assign finder_7_io_data_9 = TBEAddr_9; // @[TBE.scala 101:23]
  assign finder_7_io_data_10 = TBEAddr_10; // @[TBE.scala 101:23]
  assign finder_7_io_data_11 = TBEAddr_11; // @[TBE.scala 101:23]
  assign finder_7_io_data_12 = TBEAddr_12; // @[TBE.scala 101:23]
  assign finder_7_io_data_13 = TBEAddr_13; // @[TBE.scala 101:23]
  assign finder_7_io_data_14 = TBEAddr_14; // @[TBE.scala 101:23]
  assign finder_7_io_data_15 = TBEAddr_15; // @[TBE.scala 101:23]
  assign finder_7_io_valid_0 = TBEValid_0; // @[TBE.scala 102:24]
  assign finder_7_io_valid_1 = TBEValid_1; // @[TBE.scala 102:24]
  assign finder_7_io_valid_2 = TBEValid_2; // @[TBE.scala 102:24]
  assign finder_7_io_valid_3 = TBEValid_3; // @[TBE.scala 102:24]
  assign finder_7_io_valid_4 = TBEValid_4; // @[TBE.scala 102:24]
  assign finder_7_io_valid_5 = TBEValid_5; // @[TBE.scala 102:24]
  assign finder_7_io_valid_6 = TBEValid_6; // @[TBE.scala 102:24]
  assign finder_7_io_valid_7 = TBEValid_7; // @[TBE.scala 102:24]
  assign finder_7_io_valid_8 = TBEValid_8; // @[TBE.scala 102:24]
  assign finder_7_io_valid_9 = TBEValid_9; // @[TBE.scala 102:24]
  assign finder_7_io_valid_10 = TBEValid_10; // @[TBE.scala 102:24]
  assign finder_7_io_valid_11 = TBEValid_11; // @[TBE.scala 102:24]
  assign finder_7_io_valid_12 = TBEValid_12; // @[TBE.scala 102:24]
  assign finder_7_io_valid_13 = TBEValid_13; // @[TBE.scala 102:24]
  assign finder_7_io_valid_14 = TBEValid_14; // @[TBE.scala 102:24]
  assign finder_7_io_valid_15 = TBEValid_15; // @[TBE.scala 102:24]
  assign finder_8_io_key = io_read_bits_addr[31:0]; // @[TBE.scala 92:25]
  assign finder_8_io_data_0 = TBEAddr_0; // @[TBE.scala 93:26]
  assign finder_8_io_data_1 = TBEAddr_1; // @[TBE.scala 93:26]
  assign finder_8_io_data_2 = TBEAddr_2; // @[TBE.scala 93:26]
  assign finder_8_io_data_3 = TBEAddr_3; // @[TBE.scala 93:26]
  assign finder_8_io_data_4 = TBEAddr_4; // @[TBE.scala 93:26]
  assign finder_8_io_data_5 = TBEAddr_5; // @[TBE.scala 93:26]
  assign finder_8_io_data_6 = TBEAddr_6; // @[TBE.scala 93:26]
  assign finder_8_io_data_7 = TBEAddr_7; // @[TBE.scala 93:26]
  assign finder_8_io_data_8 = TBEAddr_8; // @[TBE.scala 93:26]
  assign finder_8_io_data_9 = TBEAddr_9; // @[TBE.scala 93:26]
  assign finder_8_io_data_10 = TBEAddr_10; // @[TBE.scala 93:26]
  assign finder_8_io_data_11 = TBEAddr_11; // @[TBE.scala 93:26]
  assign finder_8_io_data_12 = TBEAddr_12; // @[TBE.scala 93:26]
  assign finder_8_io_data_13 = TBEAddr_13; // @[TBE.scala 93:26]
  assign finder_8_io_data_14 = TBEAddr_14; // @[TBE.scala 93:26]
  assign finder_8_io_data_15 = TBEAddr_15; // @[TBE.scala 93:26]
  assign finder_8_io_valid_0 = TBEValid_0; // @[TBE.scala 94:27]
  assign finder_8_io_valid_1 = TBEValid_1; // @[TBE.scala 94:27]
  assign finder_8_io_valid_2 = TBEValid_2; // @[TBE.scala 94:27]
  assign finder_8_io_valid_3 = TBEValid_3; // @[TBE.scala 94:27]
  assign finder_8_io_valid_4 = TBEValid_4; // @[TBE.scala 94:27]
  assign finder_8_io_valid_5 = TBEValid_5; // @[TBE.scala 94:27]
  assign finder_8_io_valid_6 = TBEValid_6; // @[TBE.scala 94:27]
  assign finder_8_io_valid_7 = TBEValid_7; // @[TBE.scala 94:27]
  assign finder_8_io_valid_8 = TBEValid_8; // @[TBE.scala 94:27]
  assign finder_8_io_valid_9 = TBEValid_9; // @[TBE.scala 94:27]
  assign finder_8_io_valid_10 = TBEValid_10; // @[TBE.scala 94:27]
  assign finder_8_io_valid_11 = TBEValid_11; // @[TBE.scala 94:27]
  assign finder_8_io_valid_12 = TBEValid_12; // @[TBE.scala 94:27]
  assign finder_8_io_valid_13 = TBEValid_13; // @[TBE.scala 94:27]
  assign finder_8_io_valid_14 = TBEValid_14; // @[TBE.scala 94:27]
  assign finder_8_io_valid_15 = TBEValid_15; // @[TBE.scala 94:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  TBEMemory_0_state_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  TBEMemory_0_way = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  TBEMemory_0_fields_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  TBEMemory_1_state_state = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  TBEMemory_1_way = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  TBEMemory_1_fields_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  TBEMemory_2_state_state = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  TBEMemory_2_way = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  TBEMemory_2_fields_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  TBEMemory_3_state_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  TBEMemory_3_way = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  TBEMemory_3_fields_0 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  TBEMemory_4_state_state = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  TBEMemory_4_way = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  TBEMemory_4_fields_0 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  TBEMemory_5_state_state = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  TBEMemory_5_way = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  TBEMemory_5_fields_0 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  TBEMemory_6_state_state = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  TBEMemory_6_way = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  TBEMemory_6_fields_0 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  TBEMemory_7_state_state = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  TBEMemory_7_way = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  TBEMemory_7_fields_0 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  TBEMemory_8_state_state = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  TBEMemory_8_way = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  TBEMemory_8_fields_0 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  TBEMemory_9_state_state = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  TBEMemory_9_way = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  TBEMemory_9_fields_0 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  TBEMemory_10_state_state = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  TBEMemory_10_way = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  TBEMemory_10_fields_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  TBEMemory_11_state_state = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  TBEMemory_11_way = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  TBEMemory_11_fields_0 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  TBEMemory_12_state_state = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  TBEMemory_12_way = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  TBEMemory_12_fields_0 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  TBEMemory_13_state_state = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  TBEMemory_13_way = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  TBEMemory_13_fields_0 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  TBEMemory_14_state_state = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  TBEMemory_14_way = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  TBEMemory_14_fields_0 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  TBEMemory_15_state_state = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  TBEMemory_15_way = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  TBEMemory_15_fields_0 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  TBEValid_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  TBEValid_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  TBEValid_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  TBEValid_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  TBEValid_4 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  TBEValid_5 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  TBEValid_6 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  TBEValid_7 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  TBEValid_8 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  TBEValid_9 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  TBEValid_10 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  TBEValid_11 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  TBEValid_12 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  TBEValid_13 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  TBEValid_14 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  TBEValid_15 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  TBEAddr_0 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  TBEAddr_1 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  TBEAddr_2 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  TBEAddr_3 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  TBEAddr_4 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  TBEAddr_5 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  TBEAddr_6 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  TBEAddr_7 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  TBEAddr_8 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  TBEAddr_9 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  TBEAddr_10 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  TBEAddr_11 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  TBEAddr_12 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  TBEAddr_13 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  TBEAddr_14 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  TBEAddr_15 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  counter = _RAND_80[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      TBEMemory_0_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'h0 == idxAlloc[3:0]) begin
        TBEMemory_0_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h0 == idxAlloc[3:0]) begin
          TBEMemory_0_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEMemory_0_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEMemory_0_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEMemory_0_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEMemory_0_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEMemory_0_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEMemory_0_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEMemory_0_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h0 == idxUpdate_0[3:0]) begin
                        TBEMemory_0_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEMemory_0_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEMemory_0_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h0 == idxUpdate_0[3:0]) begin
                        TBEMemory_0_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h0 == idxAlloc[3:0]) begin
                        TBEMemory_0_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'h0 == idxUpdate_0[3:0]) begin
                        TBEMemory_0_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h0 == idxUpdate_0[3:0]) begin
                          TBEMemory_0_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEMemory_0_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEMemory_0_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h0 == idxUpdate_0[3:0]) begin
                        TBEMemory_0_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_0_state_state <= _GEN_465;
                end
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEMemory_0_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_0_state_state <= _GEN_465;
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_state_state <= 2'h0;
                  end else begin
                    TBEMemory_0_state_state <= _GEN_465;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_0_state_state <= _GEN_465;
                  end else if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_0_state_state <= _GEN_465;
                  end
                end else begin
                  TBEMemory_0_state_state <= _GEN_465;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEMemory_0_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_0_state_state <= _GEN_465;
                    end
                  end else if (_T_111) begin
                    if (4'h0 == idxUpdate_1[3:0]) begin
                      TBEMemory_0_state_state <= 2'h0;
                    end else begin
                      TBEMemory_0_state_state <= _GEN_465;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_0_state_state <= _GEN_465;
                    end else if (4'h0 == idxUpdate_1[3:0]) begin
                      TBEMemory_0_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_0_state_state <= _GEN_465;
                    end
                  end else begin
                    TBEMemory_0_state_state <= _GEN_465;
                  end
                end else if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEMemory_0_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_0_state_state <= _GEN_465;
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_state_state <= 2'h0;
                  end else begin
                    TBEMemory_0_state_state <= _GEN_465;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_0_state_state <= _GEN_465;
                  end else if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_0_state_state <= _GEN_465;
                  end
                end else begin
                  TBEMemory_0_state_state <= _GEN_465;
                end
              end else begin
                TBEMemory_0_state_state <= _GEN_979;
              end
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEMemory_0_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_0_state_state <= _GEN_979;
                end
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_state_state <= 2'h0;
                end else begin
                  TBEMemory_0_state_state <= _GEN_979;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_0_state_state <= _GEN_979;
                end else if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_0_state_state <= _GEN_979;
                end
              end else begin
                TBEMemory_0_state_state <= _GEN_979;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEMemory_0_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_0_state_state <= _GEN_979;
                  end
                end else if (_T_133) begin
                  if (4'h0 == idxUpdate_2[3:0]) begin
                    TBEMemory_0_state_state <= 2'h0;
                  end else begin
                    TBEMemory_0_state_state <= _GEN_979;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_0_state_state <= _GEN_979;
                  end else if (4'h0 == idxUpdate_2[3:0]) begin
                    TBEMemory_0_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_0_state_state <= _GEN_979;
                  end
                end else begin
                  TBEMemory_0_state_state <= _GEN_979;
                end
              end else if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEMemory_0_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_0_state_state <= _GEN_979;
                end
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_state_state <= 2'h0;
                end else begin
                  TBEMemory_0_state_state <= _GEN_979;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_0_state_state <= _GEN_979;
                end else if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_0_state_state <= _GEN_979;
                end
              end else begin
                TBEMemory_0_state_state <= _GEN_979;
              end
            end else begin
              TBEMemory_0_state_state <= _GEN_1493;
            end
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEMemory_0_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_0_state_state <= _GEN_1493;
              end
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_state_state <= 2'h0;
              end else begin
                TBEMemory_0_state_state <= _GEN_1493;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_0_state_state <= _GEN_1493;
              end else if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_0_state_state <= _GEN_1493;
              end
            end else begin
              TBEMemory_0_state_state <= _GEN_1493;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEMemory_0_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_0_state_state <= _GEN_1493;
                end
              end else if (_T_155) begin
                if (4'h0 == idxUpdate_3[3:0]) begin
                  TBEMemory_0_state_state <= 2'h0;
                end else begin
                  TBEMemory_0_state_state <= _GEN_1493;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_0_state_state <= _GEN_1493;
                end else if (4'h0 == idxUpdate_3[3:0]) begin
                  TBEMemory_0_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_0_state_state <= _GEN_1493;
                end
              end else begin
                TBEMemory_0_state_state <= _GEN_1493;
              end
            end else if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEMemory_0_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_0_state_state <= _GEN_1493;
              end
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_state_state <= 2'h0;
              end else begin
                TBEMemory_0_state_state <= _GEN_1493;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_0_state_state <= _GEN_1493;
              end else if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_0_state_state <= _GEN_1493;
              end
            end else begin
              TBEMemory_0_state_state <= _GEN_1493;
            end
          end else begin
            TBEMemory_0_state_state <= _GEN_2007;
          end
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEMemory_0_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_0_state_state <= _GEN_2007;
            end
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_state_state <= 2'h0;
            end else begin
              TBEMemory_0_state_state <= _GEN_2007;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_0_state_state <= _GEN_2007;
            end else if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_0_state_state <= _GEN_2007;
            end
          end else begin
            TBEMemory_0_state_state <= _GEN_2007;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEMemory_0_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_0_state_state <= _GEN_2007;
              end
            end else if (_T_177) begin
              if (4'h0 == idxUpdate_4[3:0]) begin
                TBEMemory_0_state_state <= 2'h0;
              end else begin
                TBEMemory_0_state_state <= _GEN_2007;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_0_state_state <= _GEN_2007;
              end else if (4'h0 == idxUpdate_4[3:0]) begin
                TBEMemory_0_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_0_state_state <= _GEN_2007;
              end
            end else begin
              TBEMemory_0_state_state <= _GEN_2007;
            end
          end else if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEMemory_0_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_0_state_state <= _GEN_2007;
            end
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_state_state <= 2'h0;
            end else begin
              TBEMemory_0_state_state <= _GEN_2007;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_0_state_state <= _GEN_2007;
            end else if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_0_state_state <= _GEN_2007;
            end
          end else begin
            TBEMemory_0_state_state <= _GEN_2007;
          end
        end else begin
          TBEMemory_0_state_state <= _GEN_2521;
        end
      end else if (_T_221) begin
        if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEMemory_0_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_0_state_state <= _GEN_2521;
          end
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_state_state <= 2'h0;
          end else begin
            TBEMemory_0_state_state <= _GEN_2521;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_0_state_state <= _GEN_2521;
          end else if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_0_state_state <= _GEN_2521;
          end
        end else begin
          TBEMemory_0_state_state <= _GEN_2521;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEMemory_0_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_0_state_state <= _GEN_2521;
            end
          end else if (_T_199) begin
            if (4'h0 == idxUpdate_5[3:0]) begin
              TBEMemory_0_state_state <= 2'h0;
            end else begin
              TBEMemory_0_state_state <= _GEN_2521;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_0_state_state <= _GEN_2521;
            end else if (4'h0 == idxUpdate_5[3:0]) begin
              TBEMemory_0_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_0_state_state <= _GEN_2521;
            end
          end else begin
            TBEMemory_0_state_state <= _GEN_2521;
          end
        end else if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEMemory_0_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_0_state_state <= _GEN_2521;
          end
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_state_state <= 2'h0;
          end else begin
            TBEMemory_0_state_state <= _GEN_2521;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_0_state_state <= _GEN_2521;
          end else if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_0_state_state <= _GEN_2521;
          end
        end else begin
          TBEMemory_0_state_state <= _GEN_2521;
        end
      end else begin
        TBEMemory_0_state_state <= _GEN_3035;
      end
    end else if (_T_243) begin
      if (4'h0 == idxUpdate_7[3:0]) begin
        TBEMemory_0_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'h0 == idxAlloc[3:0]) begin
          TBEMemory_0_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_0_state_state <= _GEN_3035;
        end
      end else if (_T_221) begin
        if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_state_state <= 2'h0;
        end else begin
          TBEMemory_0_state_state <= _GEN_3035;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_0_state_state <= _GEN_3035;
        end else if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_0_state_state <= _GEN_3035;
        end
      end else begin
        TBEMemory_0_state_state <= _GEN_3035;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEMemory_0_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_0_state_state <= _GEN_3035;
          end
        end else if (_T_221) begin
          if (4'h0 == idxUpdate_6[3:0]) begin
            TBEMemory_0_state_state <= 2'h0;
          end else begin
            TBEMemory_0_state_state <= _GEN_3035;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_0_state_state <= _GEN_3035;
          end else if (4'h0 == idxUpdate_6[3:0]) begin
            TBEMemory_0_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_0_state_state <= _GEN_3035;
          end
        end else begin
          TBEMemory_0_state_state <= _GEN_3035;
        end
      end else if (4'h0 == idxUpdate_7[3:0]) begin
        TBEMemory_0_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h0 == idxAlloc[3:0]) begin
          TBEMemory_0_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_0_state_state <= _GEN_3035;
        end
      end else if (_T_221) begin
        if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_state_state <= 2'h0;
        end else begin
          TBEMemory_0_state_state <= _GEN_3035;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_0_state_state <= _GEN_3035;
        end else if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_0_state_state <= _GEN_3035;
        end
      end else begin
        TBEMemory_0_state_state <= _GEN_3035;
      end
    end else begin
      TBEMemory_0_state_state <= _GEN_3549;
    end
    if (reset) begin
      TBEMemory_0_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'h0 == idxAlloc[3:0]) begin
        TBEMemory_0_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h0 == idxAlloc[3:0]) begin
          TBEMemory_0_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEMemory_0_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEMemory_0_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEMemory_0_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEMemory_0_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEMemory_0_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEMemory_0_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEMemory_0_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h0 == idxUpdate_0[3:0]) begin
                        TBEMemory_0_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEMemory_0_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEMemory_0_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h0 == idxUpdate_0[3:0]) begin
                        TBEMemory_0_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h0 == idxAlloc[3:0]) begin
                        TBEMemory_0_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'h0 == idxUpdate_0[3:0]) begin
                        TBEMemory_0_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h0 == idxUpdate_0[3:0]) begin
                          TBEMemory_0_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEMemory_0_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEMemory_0_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h0 == idxUpdate_0[3:0]) begin
                        TBEMemory_0_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_0_way <= _GEN_449;
                end
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEMemory_0_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_0_way <= _GEN_449;
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_way <= 3'h2;
                  end else begin
                    TBEMemory_0_way <= _GEN_449;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_0_way <= _GEN_449;
                  end else if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_0_way <= _GEN_449;
                  end
                end else begin
                  TBEMemory_0_way <= _GEN_449;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEMemory_0_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_0_way <= _GEN_449;
                    end
                  end else if (_T_111) begin
                    if (4'h0 == idxUpdate_1[3:0]) begin
                      TBEMemory_0_way <= 3'h2;
                    end else begin
                      TBEMemory_0_way <= _GEN_449;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_0_way <= _GEN_449;
                    end else if (4'h0 == idxUpdate_1[3:0]) begin
                      TBEMemory_0_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_0_way <= _GEN_449;
                    end
                  end else begin
                    TBEMemory_0_way <= _GEN_449;
                  end
                end else if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEMemory_0_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_0_way <= _GEN_449;
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_way <= 3'h2;
                  end else begin
                    TBEMemory_0_way <= _GEN_449;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_0_way <= _GEN_449;
                  end else if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_0_way <= _GEN_449;
                  end
                end else begin
                  TBEMemory_0_way <= _GEN_449;
                end
              end else begin
                TBEMemory_0_way <= _GEN_963;
              end
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEMemory_0_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_0_way <= _GEN_963;
                end
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_way <= 3'h2;
                end else begin
                  TBEMemory_0_way <= _GEN_963;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_0_way <= _GEN_963;
                end else if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_0_way <= _GEN_963;
                end
              end else begin
                TBEMemory_0_way <= _GEN_963;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEMemory_0_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_0_way <= _GEN_963;
                  end
                end else if (_T_133) begin
                  if (4'h0 == idxUpdate_2[3:0]) begin
                    TBEMemory_0_way <= 3'h2;
                  end else begin
                    TBEMemory_0_way <= _GEN_963;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_0_way <= _GEN_963;
                  end else if (4'h0 == idxUpdate_2[3:0]) begin
                    TBEMemory_0_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_0_way <= _GEN_963;
                  end
                end else begin
                  TBEMemory_0_way <= _GEN_963;
                end
              end else if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEMemory_0_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_0_way <= _GEN_963;
                end
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_way <= 3'h2;
                end else begin
                  TBEMemory_0_way <= _GEN_963;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_0_way <= _GEN_963;
                end else if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_0_way <= _GEN_963;
                end
              end else begin
                TBEMemory_0_way <= _GEN_963;
              end
            end else begin
              TBEMemory_0_way <= _GEN_1477;
            end
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEMemory_0_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_0_way <= _GEN_1477;
              end
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_way <= 3'h2;
              end else begin
                TBEMemory_0_way <= _GEN_1477;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_0_way <= _GEN_1477;
              end else if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_0_way <= _GEN_1477;
              end
            end else begin
              TBEMemory_0_way <= _GEN_1477;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEMemory_0_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_0_way <= _GEN_1477;
                end
              end else if (_T_155) begin
                if (4'h0 == idxUpdate_3[3:0]) begin
                  TBEMemory_0_way <= 3'h2;
                end else begin
                  TBEMemory_0_way <= _GEN_1477;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_0_way <= _GEN_1477;
                end else if (4'h0 == idxUpdate_3[3:0]) begin
                  TBEMemory_0_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_0_way <= _GEN_1477;
                end
              end else begin
                TBEMemory_0_way <= _GEN_1477;
              end
            end else if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEMemory_0_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_0_way <= _GEN_1477;
              end
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_way <= 3'h2;
              end else begin
                TBEMemory_0_way <= _GEN_1477;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_0_way <= _GEN_1477;
              end else if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_0_way <= _GEN_1477;
              end
            end else begin
              TBEMemory_0_way <= _GEN_1477;
            end
          end else begin
            TBEMemory_0_way <= _GEN_1991;
          end
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEMemory_0_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_0_way <= _GEN_1991;
            end
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_way <= 3'h2;
            end else begin
              TBEMemory_0_way <= _GEN_1991;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_0_way <= _GEN_1991;
            end else if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_0_way <= _GEN_1991;
            end
          end else begin
            TBEMemory_0_way <= _GEN_1991;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEMemory_0_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_0_way <= _GEN_1991;
              end
            end else if (_T_177) begin
              if (4'h0 == idxUpdate_4[3:0]) begin
                TBEMemory_0_way <= 3'h2;
              end else begin
                TBEMemory_0_way <= _GEN_1991;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_0_way <= _GEN_1991;
              end else if (4'h0 == idxUpdate_4[3:0]) begin
                TBEMemory_0_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_0_way <= _GEN_1991;
              end
            end else begin
              TBEMemory_0_way <= _GEN_1991;
            end
          end else if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEMemory_0_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_0_way <= _GEN_1991;
            end
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_way <= 3'h2;
            end else begin
              TBEMemory_0_way <= _GEN_1991;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_0_way <= _GEN_1991;
            end else if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_0_way <= _GEN_1991;
            end
          end else begin
            TBEMemory_0_way <= _GEN_1991;
          end
        end else begin
          TBEMemory_0_way <= _GEN_2505;
        end
      end else if (_T_221) begin
        if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEMemory_0_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_0_way <= _GEN_2505;
          end
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_way <= 3'h2;
          end else begin
            TBEMemory_0_way <= _GEN_2505;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_0_way <= _GEN_2505;
          end else if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_0_way <= _GEN_2505;
          end
        end else begin
          TBEMemory_0_way <= _GEN_2505;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEMemory_0_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_0_way <= _GEN_2505;
            end
          end else if (_T_199) begin
            if (4'h0 == idxUpdate_5[3:0]) begin
              TBEMemory_0_way <= 3'h2;
            end else begin
              TBEMemory_0_way <= _GEN_2505;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_0_way <= _GEN_2505;
            end else if (4'h0 == idxUpdate_5[3:0]) begin
              TBEMemory_0_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_0_way <= _GEN_2505;
            end
          end else begin
            TBEMemory_0_way <= _GEN_2505;
          end
        end else if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEMemory_0_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_0_way <= _GEN_2505;
          end
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_way <= 3'h2;
          end else begin
            TBEMemory_0_way <= _GEN_2505;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_0_way <= _GEN_2505;
          end else if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_0_way <= _GEN_2505;
          end
        end else begin
          TBEMemory_0_way <= _GEN_2505;
        end
      end else begin
        TBEMemory_0_way <= _GEN_3019;
      end
    end else if (_T_243) begin
      if (4'h0 == idxUpdate_7[3:0]) begin
        TBEMemory_0_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'h0 == idxAlloc[3:0]) begin
          TBEMemory_0_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_0_way <= _GEN_3019;
        end
      end else if (_T_221) begin
        if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_way <= 3'h2;
        end else begin
          TBEMemory_0_way <= _GEN_3019;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_0_way <= _GEN_3019;
        end else if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_0_way <= _GEN_3019;
        end
      end else begin
        TBEMemory_0_way <= _GEN_3019;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEMemory_0_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_0_way <= _GEN_3019;
          end
        end else if (_T_221) begin
          if (4'h0 == idxUpdate_6[3:0]) begin
            TBEMemory_0_way <= 3'h2;
          end else begin
            TBEMemory_0_way <= _GEN_3019;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_0_way <= _GEN_3019;
          end else if (4'h0 == idxUpdate_6[3:0]) begin
            TBEMemory_0_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_0_way <= _GEN_3019;
          end
        end else begin
          TBEMemory_0_way <= _GEN_3019;
        end
      end else if (4'h0 == idxUpdate_7[3:0]) begin
        TBEMemory_0_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h0 == idxAlloc[3:0]) begin
          TBEMemory_0_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_0_way <= _GEN_3019;
        end
      end else if (_T_221) begin
        if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_way <= 3'h2;
        end else begin
          TBEMemory_0_way <= _GEN_3019;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_0_way <= _GEN_3019;
        end else if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_0_way <= _GEN_3019;
        end
      end else begin
        TBEMemory_0_way <= _GEN_3019;
      end
    end else begin
      TBEMemory_0_way <= _GEN_3533;
    end
    if (reset) begin
      TBEMemory_0_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h0 == idxAlloc[3:0]) begin
        TBEMemory_0_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'h0 == idxAlloc[3:0]) begin
          TBEMemory_0_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEMemory_0_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEMemory_0_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEMemory_0_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEMemory_0_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEMemory_0_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEMemory_0_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEMemory_0_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h0 == idxUpdate_0[3:0]) begin
                        TBEMemory_0_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEMemory_0_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEMemory_0_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h0 == idxUpdate_0[3:0]) begin
                        TBEMemory_0_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h0 == idxUpdate_1[3:0]) begin
                      TBEMemory_0_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'h0 == idxAlloc[3:0]) begin
                        TBEMemory_0_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'h0 == idxUpdate_0[3:0]) begin
                        TBEMemory_0_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'h0 == idxUpdate_0[3:0]) begin
                          TBEMemory_0_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEMemory_0_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEMemory_0_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h0 == idxUpdate_0[3:0]) begin
                        TBEMemory_0_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_433;
                end
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEMemory_0_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_433;
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_433;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h0 == idxUpdate_1[3:0]) begin
                      TBEMemory_0_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_0_fields_0 <= _GEN_433;
                    end
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_433;
                  end
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_433;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h0 == idxUpdate_2[3:0]) begin
                    TBEMemory_0_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEMemory_0_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_0_fields_0 <= _GEN_433;
                    end
                  end else if (_T_111) begin
                    if (4'h0 == idxUpdate_1[3:0]) begin
                      TBEMemory_0_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_0_fields_0 <= _GEN_433;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'h0 == idxUpdate_1[3:0]) begin
                        TBEMemory_0_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_0_fields_0 <= _GEN_433;
                      end
                    end else begin
                      TBEMemory_0_fields_0 <= _GEN_433;
                    end
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_433;
                  end
                end else if (isAlloc_1) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEMemory_0_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_433;
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEMemory_0_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_433;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h0 == idxUpdate_1[3:0]) begin
                      TBEMemory_0_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_0_fields_0 <= _GEN_433;
                    end
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_433;
                  end
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_433;
                end
              end else begin
                TBEMemory_0_fields_0 <= _GEN_947;
              end
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEMemory_0_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_947;
                end
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_947;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h0 == idxUpdate_2[3:0]) begin
                    TBEMemory_0_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_947;
                  end
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_947;
                end
              end else begin
                TBEMemory_0_fields_0 <= _GEN_947;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h0 == idxUpdate_3[3:0]) begin
                  TBEMemory_0_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEMemory_0_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_947;
                  end
                end else if (_T_133) begin
                  if (4'h0 == idxUpdate_2[3:0]) begin
                    TBEMemory_0_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_947;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'h0 == idxUpdate_2[3:0]) begin
                      TBEMemory_0_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_0_fields_0 <= _GEN_947;
                    end
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_947;
                  end
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_947;
                end
              end else if (isAlloc_2) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEMemory_0_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_947;
                end
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEMemory_0_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_947;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h0 == idxUpdate_2[3:0]) begin
                    TBEMemory_0_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_947;
                  end
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_947;
                end
              end else begin
                TBEMemory_0_fields_0 <= _GEN_947;
              end
            end else begin
              TBEMemory_0_fields_0 <= _GEN_1461;
            end
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEMemory_0_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_0_fields_0 <= _GEN_1461;
              end
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_fields_0 <= 32'h0;
              end else begin
                TBEMemory_0_fields_0 <= _GEN_1461;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h0 == idxUpdate_3[3:0]) begin
                  TBEMemory_0_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_1461;
                end
              end else begin
                TBEMemory_0_fields_0 <= _GEN_1461;
              end
            end else begin
              TBEMemory_0_fields_0 <= _GEN_1461;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h0 == idxUpdate_4[3:0]) begin
                TBEMemory_0_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEMemory_0_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_1461;
                end
              end else if (_T_155) begin
                if (4'h0 == idxUpdate_3[3:0]) begin
                  TBEMemory_0_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_1461;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'h0 == idxUpdate_3[3:0]) begin
                    TBEMemory_0_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_0_fields_0 <= _GEN_1461;
                  end
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_1461;
                end
              end else begin
                TBEMemory_0_fields_0 <= _GEN_1461;
              end
            end else if (isAlloc_3) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEMemory_0_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_0_fields_0 <= _GEN_1461;
              end
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEMemory_0_fields_0 <= 32'h0;
              end else begin
                TBEMemory_0_fields_0 <= _GEN_1461;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h0 == idxUpdate_3[3:0]) begin
                  TBEMemory_0_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_1461;
                end
              end else begin
                TBEMemory_0_fields_0 <= _GEN_1461;
              end
            end else begin
              TBEMemory_0_fields_0 <= _GEN_1461;
            end
          end else begin
            TBEMemory_0_fields_0 <= _GEN_1975;
          end
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEMemory_0_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_0_fields_0 <= _GEN_1975;
            end
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_fields_0 <= 32'h0;
            end else begin
              TBEMemory_0_fields_0 <= _GEN_1975;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h0 == idxUpdate_4[3:0]) begin
                TBEMemory_0_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_0_fields_0 <= _GEN_1975;
              end
            end else begin
              TBEMemory_0_fields_0 <= _GEN_1975;
            end
          end else begin
            TBEMemory_0_fields_0 <= _GEN_1975;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h0 == idxUpdate_5[3:0]) begin
              TBEMemory_0_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEMemory_0_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_0_fields_0 <= _GEN_1975;
              end
            end else if (_T_177) begin
              if (4'h0 == idxUpdate_4[3:0]) begin
                TBEMemory_0_fields_0 <= 32'h0;
              end else begin
                TBEMemory_0_fields_0 <= _GEN_1975;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'h0 == idxUpdate_4[3:0]) begin
                  TBEMemory_0_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_0_fields_0 <= _GEN_1975;
                end
              end else begin
                TBEMemory_0_fields_0 <= _GEN_1975;
              end
            end else begin
              TBEMemory_0_fields_0 <= _GEN_1975;
            end
          end else if (isAlloc_4) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEMemory_0_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_0_fields_0 <= _GEN_1975;
            end
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEMemory_0_fields_0 <= 32'h0;
            end else begin
              TBEMemory_0_fields_0 <= _GEN_1975;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h0 == idxUpdate_4[3:0]) begin
                TBEMemory_0_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_0_fields_0 <= _GEN_1975;
              end
            end else begin
              TBEMemory_0_fields_0 <= _GEN_1975;
            end
          end else begin
            TBEMemory_0_fields_0 <= _GEN_1975;
          end
        end else begin
          TBEMemory_0_fields_0 <= _GEN_2489;
        end
      end else if (_T_221) begin
        if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEMemory_0_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_0_fields_0 <= _GEN_2489;
          end
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_fields_0 <= 32'h0;
          end else begin
            TBEMemory_0_fields_0 <= _GEN_2489;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h0 == idxUpdate_5[3:0]) begin
              TBEMemory_0_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_0_fields_0 <= _GEN_2489;
            end
          end else begin
            TBEMemory_0_fields_0 <= _GEN_2489;
          end
        end else begin
          TBEMemory_0_fields_0 <= _GEN_2489;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h0 == idxUpdate_6[3:0]) begin
            TBEMemory_0_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEMemory_0_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_0_fields_0 <= _GEN_2489;
            end
          end else if (_T_199) begin
            if (4'h0 == idxUpdate_5[3:0]) begin
              TBEMemory_0_fields_0 <= 32'h0;
            end else begin
              TBEMemory_0_fields_0 <= _GEN_2489;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'h0 == idxUpdate_5[3:0]) begin
                TBEMemory_0_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_0_fields_0 <= _GEN_2489;
              end
            end else begin
              TBEMemory_0_fields_0 <= _GEN_2489;
            end
          end else begin
            TBEMemory_0_fields_0 <= _GEN_2489;
          end
        end else if (isAlloc_5) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEMemory_0_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_0_fields_0 <= _GEN_2489;
          end
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEMemory_0_fields_0 <= 32'h0;
          end else begin
            TBEMemory_0_fields_0 <= _GEN_2489;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h0 == idxUpdate_5[3:0]) begin
              TBEMemory_0_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_0_fields_0 <= _GEN_2489;
            end
          end else begin
            TBEMemory_0_fields_0 <= _GEN_2489;
          end
        end else begin
          TBEMemory_0_fields_0 <= _GEN_2489;
        end
      end else begin
        TBEMemory_0_fields_0 <= _GEN_3003;
      end
    end else if (_T_243) begin
      if (4'h0 == idxUpdate_7[3:0]) begin
        TBEMemory_0_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h0 == idxAlloc[3:0]) begin
          TBEMemory_0_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_0_fields_0 <= _GEN_3003;
        end
      end else if (_T_221) begin
        if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_fields_0 <= 32'h0;
        end else begin
          TBEMemory_0_fields_0 <= _GEN_3003;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h0 == idxUpdate_6[3:0]) begin
            TBEMemory_0_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_0_fields_0 <= _GEN_3003;
          end
        end else begin
          TBEMemory_0_fields_0 <= _GEN_3003;
        end
      end else begin
        TBEMemory_0_fields_0 <= _GEN_3003;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'h0 == idxUpdate_7[3:0]) begin
          TBEMemory_0_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEMemory_0_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_0_fields_0 <= _GEN_3003;
          end
        end else if (_T_221) begin
          if (4'h0 == idxUpdate_6[3:0]) begin
            TBEMemory_0_fields_0 <= 32'h0;
          end else begin
            TBEMemory_0_fields_0 <= _GEN_3003;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'h0 == idxUpdate_6[3:0]) begin
              TBEMemory_0_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_0_fields_0 <= _GEN_3003;
            end
          end else begin
            TBEMemory_0_fields_0 <= _GEN_3003;
          end
        end else begin
          TBEMemory_0_fields_0 <= _GEN_3003;
        end
      end else if (isAlloc_6) begin
        if (4'h0 == idxAlloc[3:0]) begin
          TBEMemory_0_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_0_fields_0 <= _GEN_3003;
        end
      end else if (_T_221) begin
        if (4'h0 == idxUpdate_6[3:0]) begin
          TBEMemory_0_fields_0 <= 32'h0;
        end else begin
          TBEMemory_0_fields_0 <= _GEN_3003;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h0 == idxUpdate_6[3:0]) begin
            TBEMemory_0_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_0_fields_0 <= _GEN_3003;
          end
        end else begin
          TBEMemory_0_fields_0 <= _GEN_3003;
        end
      end else begin
        TBEMemory_0_fields_0 <= _GEN_3003;
      end
    end else begin
      TBEMemory_0_fields_0 <= _GEN_3517;
    end
    if (reset) begin
      TBEMemory_1_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'h1 == idxAlloc[3:0]) begin
        TBEMemory_1_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h1 == idxAlloc[3:0]) begin
          TBEMemory_1_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEMemory_1_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEMemory_1_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEMemory_1_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEMemory_1_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEMemory_1_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEMemory_1_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEMemory_1_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h1 == idxUpdate_0[3:0]) begin
                        TBEMemory_1_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEMemory_1_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEMemory_1_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h1 == idxUpdate_0[3:0]) begin
                        TBEMemory_1_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h1 == idxAlloc[3:0]) begin
                        TBEMemory_1_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'h1 == idxUpdate_0[3:0]) begin
                        TBEMemory_1_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h1 == idxUpdate_0[3:0]) begin
                          TBEMemory_1_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEMemory_1_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEMemory_1_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h1 == idxUpdate_0[3:0]) begin
                        TBEMemory_1_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_1_state_state <= _GEN_466;
                end
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEMemory_1_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_1_state_state <= _GEN_466;
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_state_state <= 2'h0;
                  end else begin
                    TBEMemory_1_state_state <= _GEN_466;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_1_state_state <= _GEN_466;
                  end else if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_1_state_state <= _GEN_466;
                  end
                end else begin
                  TBEMemory_1_state_state <= _GEN_466;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEMemory_1_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_1_state_state <= _GEN_466;
                    end
                  end else if (_T_111) begin
                    if (4'h1 == idxUpdate_1[3:0]) begin
                      TBEMemory_1_state_state <= 2'h0;
                    end else begin
                      TBEMemory_1_state_state <= _GEN_466;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_1_state_state <= _GEN_466;
                    end else if (4'h1 == idxUpdate_1[3:0]) begin
                      TBEMemory_1_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_1_state_state <= _GEN_466;
                    end
                  end else begin
                    TBEMemory_1_state_state <= _GEN_466;
                  end
                end else if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEMemory_1_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_1_state_state <= _GEN_466;
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_state_state <= 2'h0;
                  end else begin
                    TBEMemory_1_state_state <= _GEN_466;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_1_state_state <= _GEN_466;
                  end else if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_1_state_state <= _GEN_466;
                  end
                end else begin
                  TBEMemory_1_state_state <= _GEN_466;
                end
              end else begin
                TBEMemory_1_state_state <= _GEN_980;
              end
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEMemory_1_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_1_state_state <= _GEN_980;
                end
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_state_state <= 2'h0;
                end else begin
                  TBEMemory_1_state_state <= _GEN_980;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_1_state_state <= _GEN_980;
                end else if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_1_state_state <= _GEN_980;
                end
              end else begin
                TBEMemory_1_state_state <= _GEN_980;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEMemory_1_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_1_state_state <= _GEN_980;
                  end
                end else if (_T_133) begin
                  if (4'h1 == idxUpdate_2[3:0]) begin
                    TBEMemory_1_state_state <= 2'h0;
                  end else begin
                    TBEMemory_1_state_state <= _GEN_980;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_1_state_state <= _GEN_980;
                  end else if (4'h1 == idxUpdate_2[3:0]) begin
                    TBEMemory_1_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_1_state_state <= _GEN_980;
                  end
                end else begin
                  TBEMemory_1_state_state <= _GEN_980;
                end
              end else if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEMemory_1_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_1_state_state <= _GEN_980;
                end
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_state_state <= 2'h0;
                end else begin
                  TBEMemory_1_state_state <= _GEN_980;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_1_state_state <= _GEN_980;
                end else if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_1_state_state <= _GEN_980;
                end
              end else begin
                TBEMemory_1_state_state <= _GEN_980;
              end
            end else begin
              TBEMemory_1_state_state <= _GEN_1494;
            end
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEMemory_1_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_1_state_state <= _GEN_1494;
              end
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_state_state <= 2'h0;
              end else begin
                TBEMemory_1_state_state <= _GEN_1494;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_1_state_state <= _GEN_1494;
              end else if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_1_state_state <= _GEN_1494;
              end
            end else begin
              TBEMemory_1_state_state <= _GEN_1494;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEMemory_1_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_1_state_state <= _GEN_1494;
                end
              end else if (_T_155) begin
                if (4'h1 == idxUpdate_3[3:0]) begin
                  TBEMemory_1_state_state <= 2'h0;
                end else begin
                  TBEMemory_1_state_state <= _GEN_1494;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_1_state_state <= _GEN_1494;
                end else if (4'h1 == idxUpdate_3[3:0]) begin
                  TBEMemory_1_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_1_state_state <= _GEN_1494;
                end
              end else begin
                TBEMemory_1_state_state <= _GEN_1494;
              end
            end else if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEMemory_1_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_1_state_state <= _GEN_1494;
              end
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_state_state <= 2'h0;
              end else begin
                TBEMemory_1_state_state <= _GEN_1494;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_1_state_state <= _GEN_1494;
              end else if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_1_state_state <= _GEN_1494;
              end
            end else begin
              TBEMemory_1_state_state <= _GEN_1494;
            end
          end else begin
            TBEMemory_1_state_state <= _GEN_2008;
          end
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEMemory_1_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_1_state_state <= _GEN_2008;
            end
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_state_state <= 2'h0;
            end else begin
              TBEMemory_1_state_state <= _GEN_2008;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_1_state_state <= _GEN_2008;
            end else if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_1_state_state <= _GEN_2008;
            end
          end else begin
            TBEMemory_1_state_state <= _GEN_2008;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEMemory_1_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_1_state_state <= _GEN_2008;
              end
            end else if (_T_177) begin
              if (4'h1 == idxUpdate_4[3:0]) begin
                TBEMemory_1_state_state <= 2'h0;
              end else begin
                TBEMemory_1_state_state <= _GEN_2008;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_1_state_state <= _GEN_2008;
              end else if (4'h1 == idxUpdate_4[3:0]) begin
                TBEMemory_1_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_1_state_state <= _GEN_2008;
              end
            end else begin
              TBEMemory_1_state_state <= _GEN_2008;
            end
          end else if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEMemory_1_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_1_state_state <= _GEN_2008;
            end
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_state_state <= 2'h0;
            end else begin
              TBEMemory_1_state_state <= _GEN_2008;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_1_state_state <= _GEN_2008;
            end else if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_1_state_state <= _GEN_2008;
            end
          end else begin
            TBEMemory_1_state_state <= _GEN_2008;
          end
        end else begin
          TBEMemory_1_state_state <= _GEN_2522;
        end
      end else if (_T_221) begin
        if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEMemory_1_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_1_state_state <= _GEN_2522;
          end
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_state_state <= 2'h0;
          end else begin
            TBEMemory_1_state_state <= _GEN_2522;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_1_state_state <= _GEN_2522;
          end else if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_1_state_state <= _GEN_2522;
          end
        end else begin
          TBEMemory_1_state_state <= _GEN_2522;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEMemory_1_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_1_state_state <= _GEN_2522;
            end
          end else if (_T_199) begin
            if (4'h1 == idxUpdate_5[3:0]) begin
              TBEMemory_1_state_state <= 2'h0;
            end else begin
              TBEMemory_1_state_state <= _GEN_2522;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_1_state_state <= _GEN_2522;
            end else if (4'h1 == idxUpdate_5[3:0]) begin
              TBEMemory_1_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_1_state_state <= _GEN_2522;
            end
          end else begin
            TBEMemory_1_state_state <= _GEN_2522;
          end
        end else if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEMemory_1_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_1_state_state <= _GEN_2522;
          end
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_state_state <= 2'h0;
          end else begin
            TBEMemory_1_state_state <= _GEN_2522;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_1_state_state <= _GEN_2522;
          end else if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_1_state_state <= _GEN_2522;
          end
        end else begin
          TBEMemory_1_state_state <= _GEN_2522;
        end
      end else begin
        TBEMemory_1_state_state <= _GEN_3036;
      end
    end else if (_T_243) begin
      if (4'h1 == idxUpdate_7[3:0]) begin
        TBEMemory_1_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'h1 == idxAlloc[3:0]) begin
          TBEMemory_1_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_1_state_state <= _GEN_3036;
        end
      end else if (_T_221) begin
        if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_state_state <= 2'h0;
        end else begin
          TBEMemory_1_state_state <= _GEN_3036;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_1_state_state <= _GEN_3036;
        end else if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_1_state_state <= _GEN_3036;
        end
      end else begin
        TBEMemory_1_state_state <= _GEN_3036;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEMemory_1_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_1_state_state <= _GEN_3036;
          end
        end else if (_T_221) begin
          if (4'h1 == idxUpdate_6[3:0]) begin
            TBEMemory_1_state_state <= 2'h0;
          end else begin
            TBEMemory_1_state_state <= _GEN_3036;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_1_state_state <= _GEN_3036;
          end else if (4'h1 == idxUpdate_6[3:0]) begin
            TBEMemory_1_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_1_state_state <= _GEN_3036;
          end
        end else begin
          TBEMemory_1_state_state <= _GEN_3036;
        end
      end else if (4'h1 == idxUpdate_7[3:0]) begin
        TBEMemory_1_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h1 == idxAlloc[3:0]) begin
          TBEMemory_1_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_1_state_state <= _GEN_3036;
        end
      end else if (_T_221) begin
        if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_state_state <= 2'h0;
        end else begin
          TBEMemory_1_state_state <= _GEN_3036;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_1_state_state <= _GEN_3036;
        end else if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_1_state_state <= _GEN_3036;
        end
      end else begin
        TBEMemory_1_state_state <= _GEN_3036;
      end
    end else begin
      TBEMemory_1_state_state <= _GEN_3550;
    end
    if (reset) begin
      TBEMemory_1_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'h1 == idxAlloc[3:0]) begin
        TBEMemory_1_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h1 == idxAlloc[3:0]) begin
          TBEMemory_1_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEMemory_1_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEMemory_1_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEMemory_1_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEMemory_1_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEMemory_1_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEMemory_1_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEMemory_1_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h1 == idxUpdate_0[3:0]) begin
                        TBEMemory_1_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEMemory_1_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEMemory_1_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h1 == idxUpdate_0[3:0]) begin
                        TBEMemory_1_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h1 == idxAlloc[3:0]) begin
                        TBEMemory_1_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'h1 == idxUpdate_0[3:0]) begin
                        TBEMemory_1_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h1 == idxUpdate_0[3:0]) begin
                          TBEMemory_1_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEMemory_1_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEMemory_1_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h1 == idxUpdate_0[3:0]) begin
                        TBEMemory_1_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_1_way <= _GEN_450;
                end
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEMemory_1_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_1_way <= _GEN_450;
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_way <= 3'h2;
                  end else begin
                    TBEMemory_1_way <= _GEN_450;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_1_way <= _GEN_450;
                  end else if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_1_way <= _GEN_450;
                  end
                end else begin
                  TBEMemory_1_way <= _GEN_450;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEMemory_1_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_1_way <= _GEN_450;
                    end
                  end else if (_T_111) begin
                    if (4'h1 == idxUpdate_1[3:0]) begin
                      TBEMemory_1_way <= 3'h2;
                    end else begin
                      TBEMemory_1_way <= _GEN_450;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_1_way <= _GEN_450;
                    end else if (4'h1 == idxUpdate_1[3:0]) begin
                      TBEMemory_1_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_1_way <= _GEN_450;
                    end
                  end else begin
                    TBEMemory_1_way <= _GEN_450;
                  end
                end else if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEMemory_1_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_1_way <= _GEN_450;
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_way <= 3'h2;
                  end else begin
                    TBEMemory_1_way <= _GEN_450;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_1_way <= _GEN_450;
                  end else if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_1_way <= _GEN_450;
                  end
                end else begin
                  TBEMemory_1_way <= _GEN_450;
                end
              end else begin
                TBEMemory_1_way <= _GEN_964;
              end
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEMemory_1_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_1_way <= _GEN_964;
                end
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_way <= 3'h2;
                end else begin
                  TBEMemory_1_way <= _GEN_964;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_1_way <= _GEN_964;
                end else if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_1_way <= _GEN_964;
                end
              end else begin
                TBEMemory_1_way <= _GEN_964;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEMemory_1_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_1_way <= _GEN_964;
                  end
                end else if (_T_133) begin
                  if (4'h1 == idxUpdate_2[3:0]) begin
                    TBEMemory_1_way <= 3'h2;
                  end else begin
                    TBEMemory_1_way <= _GEN_964;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_1_way <= _GEN_964;
                  end else if (4'h1 == idxUpdate_2[3:0]) begin
                    TBEMemory_1_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_1_way <= _GEN_964;
                  end
                end else begin
                  TBEMemory_1_way <= _GEN_964;
                end
              end else if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEMemory_1_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_1_way <= _GEN_964;
                end
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_way <= 3'h2;
                end else begin
                  TBEMemory_1_way <= _GEN_964;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_1_way <= _GEN_964;
                end else if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_1_way <= _GEN_964;
                end
              end else begin
                TBEMemory_1_way <= _GEN_964;
              end
            end else begin
              TBEMemory_1_way <= _GEN_1478;
            end
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEMemory_1_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_1_way <= _GEN_1478;
              end
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_way <= 3'h2;
              end else begin
                TBEMemory_1_way <= _GEN_1478;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_1_way <= _GEN_1478;
              end else if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_1_way <= _GEN_1478;
              end
            end else begin
              TBEMemory_1_way <= _GEN_1478;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEMemory_1_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_1_way <= _GEN_1478;
                end
              end else if (_T_155) begin
                if (4'h1 == idxUpdate_3[3:0]) begin
                  TBEMemory_1_way <= 3'h2;
                end else begin
                  TBEMemory_1_way <= _GEN_1478;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_1_way <= _GEN_1478;
                end else if (4'h1 == idxUpdate_3[3:0]) begin
                  TBEMemory_1_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_1_way <= _GEN_1478;
                end
              end else begin
                TBEMemory_1_way <= _GEN_1478;
              end
            end else if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEMemory_1_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_1_way <= _GEN_1478;
              end
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_way <= 3'h2;
              end else begin
                TBEMemory_1_way <= _GEN_1478;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_1_way <= _GEN_1478;
              end else if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_1_way <= _GEN_1478;
              end
            end else begin
              TBEMemory_1_way <= _GEN_1478;
            end
          end else begin
            TBEMemory_1_way <= _GEN_1992;
          end
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEMemory_1_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_1_way <= _GEN_1992;
            end
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_way <= 3'h2;
            end else begin
              TBEMemory_1_way <= _GEN_1992;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_1_way <= _GEN_1992;
            end else if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_1_way <= _GEN_1992;
            end
          end else begin
            TBEMemory_1_way <= _GEN_1992;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEMemory_1_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_1_way <= _GEN_1992;
              end
            end else if (_T_177) begin
              if (4'h1 == idxUpdate_4[3:0]) begin
                TBEMemory_1_way <= 3'h2;
              end else begin
                TBEMemory_1_way <= _GEN_1992;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_1_way <= _GEN_1992;
              end else if (4'h1 == idxUpdate_4[3:0]) begin
                TBEMemory_1_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_1_way <= _GEN_1992;
              end
            end else begin
              TBEMemory_1_way <= _GEN_1992;
            end
          end else if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEMemory_1_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_1_way <= _GEN_1992;
            end
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_way <= 3'h2;
            end else begin
              TBEMemory_1_way <= _GEN_1992;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_1_way <= _GEN_1992;
            end else if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_1_way <= _GEN_1992;
            end
          end else begin
            TBEMemory_1_way <= _GEN_1992;
          end
        end else begin
          TBEMemory_1_way <= _GEN_2506;
        end
      end else if (_T_221) begin
        if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEMemory_1_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_1_way <= _GEN_2506;
          end
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_way <= 3'h2;
          end else begin
            TBEMemory_1_way <= _GEN_2506;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_1_way <= _GEN_2506;
          end else if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_1_way <= _GEN_2506;
          end
        end else begin
          TBEMemory_1_way <= _GEN_2506;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEMemory_1_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_1_way <= _GEN_2506;
            end
          end else if (_T_199) begin
            if (4'h1 == idxUpdate_5[3:0]) begin
              TBEMemory_1_way <= 3'h2;
            end else begin
              TBEMemory_1_way <= _GEN_2506;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_1_way <= _GEN_2506;
            end else if (4'h1 == idxUpdate_5[3:0]) begin
              TBEMemory_1_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_1_way <= _GEN_2506;
            end
          end else begin
            TBEMemory_1_way <= _GEN_2506;
          end
        end else if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEMemory_1_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_1_way <= _GEN_2506;
          end
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_way <= 3'h2;
          end else begin
            TBEMemory_1_way <= _GEN_2506;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_1_way <= _GEN_2506;
          end else if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_1_way <= _GEN_2506;
          end
        end else begin
          TBEMemory_1_way <= _GEN_2506;
        end
      end else begin
        TBEMemory_1_way <= _GEN_3020;
      end
    end else if (_T_243) begin
      if (4'h1 == idxUpdate_7[3:0]) begin
        TBEMemory_1_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'h1 == idxAlloc[3:0]) begin
          TBEMemory_1_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_1_way <= _GEN_3020;
        end
      end else if (_T_221) begin
        if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_way <= 3'h2;
        end else begin
          TBEMemory_1_way <= _GEN_3020;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_1_way <= _GEN_3020;
        end else if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_1_way <= _GEN_3020;
        end
      end else begin
        TBEMemory_1_way <= _GEN_3020;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEMemory_1_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_1_way <= _GEN_3020;
          end
        end else if (_T_221) begin
          if (4'h1 == idxUpdate_6[3:0]) begin
            TBEMemory_1_way <= 3'h2;
          end else begin
            TBEMemory_1_way <= _GEN_3020;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_1_way <= _GEN_3020;
          end else if (4'h1 == idxUpdate_6[3:0]) begin
            TBEMemory_1_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_1_way <= _GEN_3020;
          end
        end else begin
          TBEMemory_1_way <= _GEN_3020;
        end
      end else if (4'h1 == idxUpdate_7[3:0]) begin
        TBEMemory_1_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h1 == idxAlloc[3:0]) begin
          TBEMemory_1_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_1_way <= _GEN_3020;
        end
      end else if (_T_221) begin
        if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_way <= 3'h2;
        end else begin
          TBEMemory_1_way <= _GEN_3020;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_1_way <= _GEN_3020;
        end else if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_1_way <= _GEN_3020;
        end
      end else begin
        TBEMemory_1_way <= _GEN_3020;
      end
    end else begin
      TBEMemory_1_way <= _GEN_3534;
    end
    if (reset) begin
      TBEMemory_1_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h1 == idxAlloc[3:0]) begin
        TBEMemory_1_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'h1 == idxAlloc[3:0]) begin
          TBEMemory_1_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEMemory_1_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEMemory_1_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEMemory_1_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEMemory_1_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEMemory_1_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEMemory_1_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEMemory_1_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h1 == idxUpdate_0[3:0]) begin
                        TBEMemory_1_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEMemory_1_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEMemory_1_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h1 == idxUpdate_0[3:0]) begin
                        TBEMemory_1_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h1 == idxUpdate_1[3:0]) begin
                      TBEMemory_1_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'h1 == idxAlloc[3:0]) begin
                        TBEMemory_1_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'h1 == idxUpdate_0[3:0]) begin
                        TBEMemory_1_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'h1 == idxUpdate_0[3:0]) begin
                          TBEMemory_1_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEMemory_1_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEMemory_1_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h1 == idxUpdate_0[3:0]) begin
                        TBEMemory_1_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_434;
                end
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEMemory_1_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_434;
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_434;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h1 == idxUpdate_1[3:0]) begin
                      TBEMemory_1_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_1_fields_0 <= _GEN_434;
                    end
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_434;
                  end
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_434;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h1 == idxUpdate_2[3:0]) begin
                    TBEMemory_1_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEMemory_1_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_1_fields_0 <= _GEN_434;
                    end
                  end else if (_T_111) begin
                    if (4'h1 == idxUpdate_1[3:0]) begin
                      TBEMemory_1_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_1_fields_0 <= _GEN_434;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'h1 == idxUpdate_1[3:0]) begin
                        TBEMemory_1_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_1_fields_0 <= _GEN_434;
                      end
                    end else begin
                      TBEMemory_1_fields_0 <= _GEN_434;
                    end
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_434;
                  end
                end else if (isAlloc_1) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEMemory_1_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_434;
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEMemory_1_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_434;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h1 == idxUpdate_1[3:0]) begin
                      TBEMemory_1_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_1_fields_0 <= _GEN_434;
                    end
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_434;
                  end
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_434;
                end
              end else begin
                TBEMemory_1_fields_0 <= _GEN_948;
              end
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEMemory_1_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_948;
                end
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_948;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h1 == idxUpdate_2[3:0]) begin
                    TBEMemory_1_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_948;
                  end
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_948;
                end
              end else begin
                TBEMemory_1_fields_0 <= _GEN_948;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h1 == idxUpdate_3[3:0]) begin
                  TBEMemory_1_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEMemory_1_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_948;
                  end
                end else if (_T_133) begin
                  if (4'h1 == idxUpdate_2[3:0]) begin
                    TBEMemory_1_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_948;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'h1 == idxUpdate_2[3:0]) begin
                      TBEMemory_1_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_1_fields_0 <= _GEN_948;
                    end
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_948;
                  end
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_948;
                end
              end else if (isAlloc_2) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEMemory_1_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_948;
                end
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEMemory_1_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_948;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h1 == idxUpdate_2[3:0]) begin
                    TBEMemory_1_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_948;
                  end
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_948;
                end
              end else begin
                TBEMemory_1_fields_0 <= _GEN_948;
              end
            end else begin
              TBEMemory_1_fields_0 <= _GEN_1462;
            end
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEMemory_1_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_1_fields_0 <= _GEN_1462;
              end
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_fields_0 <= 32'h0;
              end else begin
                TBEMemory_1_fields_0 <= _GEN_1462;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h1 == idxUpdate_3[3:0]) begin
                  TBEMemory_1_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_1462;
                end
              end else begin
                TBEMemory_1_fields_0 <= _GEN_1462;
              end
            end else begin
              TBEMemory_1_fields_0 <= _GEN_1462;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h1 == idxUpdate_4[3:0]) begin
                TBEMemory_1_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEMemory_1_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_1462;
                end
              end else if (_T_155) begin
                if (4'h1 == idxUpdate_3[3:0]) begin
                  TBEMemory_1_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_1462;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'h1 == idxUpdate_3[3:0]) begin
                    TBEMemory_1_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_1_fields_0 <= _GEN_1462;
                  end
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_1462;
                end
              end else begin
                TBEMemory_1_fields_0 <= _GEN_1462;
              end
            end else if (isAlloc_3) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEMemory_1_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_1_fields_0 <= _GEN_1462;
              end
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEMemory_1_fields_0 <= 32'h0;
              end else begin
                TBEMemory_1_fields_0 <= _GEN_1462;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h1 == idxUpdate_3[3:0]) begin
                  TBEMemory_1_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_1462;
                end
              end else begin
                TBEMemory_1_fields_0 <= _GEN_1462;
              end
            end else begin
              TBEMemory_1_fields_0 <= _GEN_1462;
            end
          end else begin
            TBEMemory_1_fields_0 <= _GEN_1976;
          end
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEMemory_1_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_1_fields_0 <= _GEN_1976;
            end
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_fields_0 <= 32'h0;
            end else begin
              TBEMemory_1_fields_0 <= _GEN_1976;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h1 == idxUpdate_4[3:0]) begin
                TBEMemory_1_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_1_fields_0 <= _GEN_1976;
              end
            end else begin
              TBEMemory_1_fields_0 <= _GEN_1976;
            end
          end else begin
            TBEMemory_1_fields_0 <= _GEN_1976;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h1 == idxUpdate_5[3:0]) begin
              TBEMemory_1_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEMemory_1_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_1_fields_0 <= _GEN_1976;
              end
            end else if (_T_177) begin
              if (4'h1 == idxUpdate_4[3:0]) begin
                TBEMemory_1_fields_0 <= 32'h0;
              end else begin
                TBEMemory_1_fields_0 <= _GEN_1976;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'h1 == idxUpdate_4[3:0]) begin
                  TBEMemory_1_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_1_fields_0 <= _GEN_1976;
                end
              end else begin
                TBEMemory_1_fields_0 <= _GEN_1976;
              end
            end else begin
              TBEMemory_1_fields_0 <= _GEN_1976;
            end
          end else if (isAlloc_4) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEMemory_1_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_1_fields_0 <= _GEN_1976;
            end
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEMemory_1_fields_0 <= 32'h0;
            end else begin
              TBEMemory_1_fields_0 <= _GEN_1976;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h1 == idxUpdate_4[3:0]) begin
                TBEMemory_1_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_1_fields_0 <= _GEN_1976;
              end
            end else begin
              TBEMemory_1_fields_0 <= _GEN_1976;
            end
          end else begin
            TBEMemory_1_fields_0 <= _GEN_1976;
          end
        end else begin
          TBEMemory_1_fields_0 <= _GEN_2490;
        end
      end else if (_T_221) begin
        if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEMemory_1_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_1_fields_0 <= _GEN_2490;
          end
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_fields_0 <= 32'h0;
          end else begin
            TBEMemory_1_fields_0 <= _GEN_2490;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h1 == idxUpdate_5[3:0]) begin
              TBEMemory_1_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_1_fields_0 <= _GEN_2490;
            end
          end else begin
            TBEMemory_1_fields_0 <= _GEN_2490;
          end
        end else begin
          TBEMemory_1_fields_0 <= _GEN_2490;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h1 == idxUpdate_6[3:0]) begin
            TBEMemory_1_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEMemory_1_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_1_fields_0 <= _GEN_2490;
            end
          end else if (_T_199) begin
            if (4'h1 == idxUpdate_5[3:0]) begin
              TBEMemory_1_fields_0 <= 32'h0;
            end else begin
              TBEMemory_1_fields_0 <= _GEN_2490;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'h1 == idxUpdate_5[3:0]) begin
                TBEMemory_1_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_1_fields_0 <= _GEN_2490;
              end
            end else begin
              TBEMemory_1_fields_0 <= _GEN_2490;
            end
          end else begin
            TBEMemory_1_fields_0 <= _GEN_2490;
          end
        end else if (isAlloc_5) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEMemory_1_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_1_fields_0 <= _GEN_2490;
          end
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEMemory_1_fields_0 <= 32'h0;
          end else begin
            TBEMemory_1_fields_0 <= _GEN_2490;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h1 == idxUpdate_5[3:0]) begin
              TBEMemory_1_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_1_fields_0 <= _GEN_2490;
            end
          end else begin
            TBEMemory_1_fields_0 <= _GEN_2490;
          end
        end else begin
          TBEMemory_1_fields_0 <= _GEN_2490;
        end
      end else begin
        TBEMemory_1_fields_0 <= _GEN_3004;
      end
    end else if (_T_243) begin
      if (4'h1 == idxUpdate_7[3:0]) begin
        TBEMemory_1_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h1 == idxAlloc[3:0]) begin
          TBEMemory_1_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_1_fields_0 <= _GEN_3004;
        end
      end else if (_T_221) begin
        if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_fields_0 <= 32'h0;
        end else begin
          TBEMemory_1_fields_0 <= _GEN_3004;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h1 == idxUpdate_6[3:0]) begin
            TBEMemory_1_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_1_fields_0 <= _GEN_3004;
          end
        end else begin
          TBEMemory_1_fields_0 <= _GEN_3004;
        end
      end else begin
        TBEMemory_1_fields_0 <= _GEN_3004;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'h1 == idxUpdate_7[3:0]) begin
          TBEMemory_1_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEMemory_1_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_1_fields_0 <= _GEN_3004;
          end
        end else if (_T_221) begin
          if (4'h1 == idxUpdate_6[3:0]) begin
            TBEMemory_1_fields_0 <= 32'h0;
          end else begin
            TBEMemory_1_fields_0 <= _GEN_3004;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'h1 == idxUpdate_6[3:0]) begin
              TBEMemory_1_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_1_fields_0 <= _GEN_3004;
            end
          end else begin
            TBEMemory_1_fields_0 <= _GEN_3004;
          end
        end else begin
          TBEMemory_1_fields_0 <= _GEN_3004;
        end
      end else if (isAlloc_6) begin
        if (4'h1 == idxAlloc[3:0]) begin
          TBEMemory_1_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_1_fields_0 <= _GEN_3004;
        end
      end else if (_T_221) begin
        if (4'h1 == idxUpdate_6[3:0]) begin
          TBEMemory_1_fields_0 <= 32'h0;
        end else begin
          TBEMemory_1_fields_0 <= _GEN_3004;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h1 == idxUpdate_6[3:0]) begin
            TBEMemory_1_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_1_fields_0 <= _GEN_3004;
          end
        end else begin
          TBEMemory_1_fields_0 <= _GEN_3004;
        end
      end else begin
        TBEMemory_1_fields_0 <= _GEN_3004;
      end
    end else begin
      TBEMemory_1_fields_0 <= _GEN_3518;
    end
    if (reset) begin
      TBEMemory_2_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'h2 == idxAlloc[3:0]) begin
        TBEMemory_2_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h2 == idxAlloc[3:0]) begin
          TBEMemory_2_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEMemory_2_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEMemory_2_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEMemory_2_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEMemory_2_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEMemory_2_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEMemory_2_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEMemory_2_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h2 == idxUpdate_0[3:0]) begin
                        TBEMemory_2_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEMemory_2_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEMemory_2_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h2 == idxUpdate_0[3:0]) begin
                        TBEMemory_2_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h2 == idxAlloc[3:0]) begin
                        TBEMemory_2_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'h2 == idxUpdate_0[3:0]) begin
                        TBEMemory_2_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h2 == idxUpdate_0[3:0]) begin
                          TBEMemory_2_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEMemory_2_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEMemory_2_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h2 == idxUpdate_0[3:0]) begin
                        TBEMemory_2_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_2_state_state <= _GEN_467;
                end
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEMemory_2_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_2_state_state <= _GEN_467;
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_state_state <= 2'h0;
                  end else begin
                    TBEMemory_2_state_state <= _GEN_467;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_2_state_state <= _GEN_467;
                  end else if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_2_state_state <= _GEN_467;
                  end
                end else begin
                  TBEMemory_2_state_state <= _GEN_467;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEMemory_2_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_2_state_state <= _GEN_467;
                    end
                  end else if (_T_111) begin
                    if (4'h2 == idxUpdate_1[3:0]) begin
                      TBEMemory_2_state_state <= 2'h0;
                    end else begin
                      TBEMemory_2_state_state <= _GEN_467;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_2_state_state <= _GEN_467;
                    end else if (4'h2 == idxUpdate_1[3:0]) begin
                      TBEMemory_2_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_2_state_state <= _GEN_467;
                    end
                  end else begin
                    TBEMemory_2_state_state <= _GEN_467;
                  end
                end else if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEMemory_2_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_2_state_state <= _GEN_467;
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_state_state <= 2'h0;
                  end else begin
                    TBEMemory_2_state_state <= _GEN_467;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_2_state_state <= _GEN_467;
                  end else if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_2_state_state <= _GEN_467;
                  end
                end else begin
                  TBEMemory_2_state_state <= _GEN_467;
                end
              end else begin
                TBEMemory_2_state_state <= _GEN_981;
              end
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEMemory_2_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_2_state_state <= _GEN_981;
                end
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_state_state <= 2'h0;
                end else begin
                  TBEMemory_2_state_state <= _GEN_981;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_2_state_state <= _GEN_981;
                end else if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_2_state_state <= _GEN_981;
                end
              end else begin
                TBEMemory_2_state_state <= _GEN_981;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEMemory_2_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_2_state_state <= _GEN_981;
                  end
                end else if (_T_133) begin
                  if (4'h2 == idxUpdate_2[3:0]) begin
                    TBEMemory_2_state_state <= 2'h0;
                  end else begin
                    TBEMemory_2_state_state <= _GEN_981;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_2_state_state <= _GEN_981;
                  end else if (4'h2 == idxUpdate_2[3:0]) begin
                    TBEMemory_2_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_2_state_state <= _GEN_981;
                  end
                end else begin
                  TBEMemory_2_state_state <= _GEN_981;
                end
              end else if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEMemory_2_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_2_state_state <= _GEN_981;
                end
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_state_state <= 2'h0;
                end else begin
                  TBEMemory_2_state_state <= _GEN_981;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_2_state_state <= _GEN_981;
                end else if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_2_state_state <= _GEN_981;
                end
              end else begin
                TBEMemory_2_state_state <= _GEN_981;
              end
            end else begin
              TBEMemory_2_state_state <= _GEN_1495;
            end
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEMemory_2_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_2_state_state <= _GEN_1495;
              end
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_state_state <= 2'h0;
              end else begin
                TBEMemory_2_state_state <= _GEN_1495;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_2_state_state <= _GEN_1495;
              end else if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_2_state_state <= _GEN_1495;
              end
            end else begin
              TBEMemory_2_state_state <= _GEN_1495;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEMemory_2_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_2_state_state <= _GEN_1495;
                end
              end else if (_T_155) begin
                if (4'h2 == idxUpdate_3[3:0]) begin
                  TBEMemory_2_state_state <= 2'h0;
                end else begin
                  TBEMemory_2_state_state <= _GEN_1495;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_2_state_state <= _GEN_1495;
                end else if (4'h2 == idxUpdate_3[3:0]) begin
                  TBEMemory_2_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_2_state_state <= _GEN_1495;
                end
              end else begin
                TBEMemory_2_state_state <= _GEN_1495;
              end
            end else if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEMemory_2_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_2_state_state <= _GEN_1495;
              end
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_state_state <= 2'h0;
              end else begin
                TBEMemory_2_state_state <= _GEN_1495;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_2_state_state <= _GEN_1495;
              end else if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_2_state_state <= _GEN_1495;
              end
            end else begin
              TBEMemory_2_state_state <= _GEN_1495;
            end
          end else begin
            TBEMemory_2_state_state <= _GEN_2009;
          end
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEMemory_2_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_2_state_state <= _GEN_2009;
            end
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_state_state <= 2'h0;
            end else begin
              TBEMemory_2_state_state <= _GEN_2009;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_2_state_state <= _GEN_2009;
            end else if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_2_state_state <= _GEN_2009;
            end
          end else begin
            TBEMemory_2_state_state <= _GEN_2009;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEMemory_2_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_2_state_state <= _GEN_2009;
              end
            end else if (_T_177) begin
              if (4'h2 == idxUpdate_4[3:0]) begin
                TBEMemory_2_state_state <= 2'h0;
              end else begin
                TBEMemory_2_state_state <= _GEN_2009;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_2_state_state <= _GEN_2009;
              end else if (4'h2 == idxUpdate_4[3:0]) begin
                TBEMemory_2_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_2_state_state <= _GEN_2009;
              end
            end else begin
              TBEMemory_2_state_state <= _GEN_2009;
            end
          end else if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEMemory_2_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_2_state_state <= _GEN_2009;
            end
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_state_state <= 2'h0;
            end else begin
              TBEMemory_2_state_state <= _GEN_2009;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_2_state_state <= _GEN_2009;
            end else if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_2_state_state <= _GEN_2009;
            end
          end else begin
            TBEMemory_2_state_state <= _GEN_2009;
          end
        end else begin
          TBEMemory_2_state_state <= _GEN_2523;
        end
      end else if (_T_221) begin
        if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEMemory_2_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_2_state_state <= _GEN_2523;
          end
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_state_state <= 2'h0;
          end else begin
            TBEMemory_2_state_state <= _GEN_2523;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_2_state_state <= _GEN_2523;
          end else if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_2_state_state <= _GEN_2523;
          end
        end else begin
          TBEMemory_2_state_state <= _GEN_2523;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEMemory_2_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_2_state_state <= _GEN_2523;
            end
          end else if (_T_199) begin
            if (4'h2 == idxUpdate_5[3:0]) begin
              TBEMemory_2_state_state <= 2'h0;
            end else begin
              TBEMemory_2_state_state <= _GEN_2523;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_2_state_state <= _GEN_2523;
            end else if (4'h2 == idxUpdate_5[3:0]) begin
              TBEMemory_2_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_2_state_state <= _GEN_2523;
            end
          end else begin
            TBEMemory_2_state_state <= _GEN_2523;
          end
        end else if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEMemory_2_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_2_state_state <= _GEN_2523;
          end
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_state_state <= 2'h0;
          end else begin
            TBEMemory_2_state_state <= _GEN_2523;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_2_state_state <= _GEN_2523;
          end else if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_2_state_state <= _GEN_2523;
          end
        end else begin
          TBEMemory_2_state_state <= _GEN_2523;
        end
      end else begin
        TBEMemory_2_state_state <= _GEN_3037;
      end
    end else if (_T_243) begin
      if (4'h2 == idxUpdate_7[3:0]) begin
        TBEMemory_2_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'h2 == idxAlloc[3:0]) begin
          TBEMemory_2_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_2_state_state <= _GEN_3037;
        end
      end else if (_T_221) begin
        if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_state_state <= 2'h0;
        end else begin
          TBEMemory_2_state_state <= _GEN_3037;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_2_state_state <= _GEN_3037;
        end else if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_2_state_state <= _GEN_3037;
        end
      end else begin
        TBEMemory_2_state_state <= _GEN_3037;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEMemory_2_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_2_state_state <= _GEN_3037;
          end
        end else if (_T_221) begin
          if (4'h2 == idxUpdate_6[3:0]) begin
            TBEMemory_2_state_state <= 2'h0;
          end else begin
            TBEMemory_2_state_state <= _GEN_3037;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_2_state_state <= _GEN_3037;
          end else if (4'h2 == idxUpdate_6[3:0]) begin
            TBEMemory_2_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_2_state_state <= _GEN_3037;
          end
        end else begin
          TBEMemory_2_state_state <= _GEN_3037;
        end
      end else if (4'h2 == idxUpdate_7[3:0]) begin
        TBEMemory_2_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h2 == idxAlloc[3:0]) begin
          TBEMemory_2_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_2_state_state <= _GEN_3037;
        end
      end else if (_T_221) begin
        if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_state_state <= 2'h0;
        end else begin
          TBEMemory_2_state_state <= _GEN_3037;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_2_state_state <= _GEN_3037;
        end else if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_2_state_state <= _GEN_3037;
        end
      end else begin
        TBEMemory_2_state_state <= _GEN_3037;
      end
    end else begin
      TBEMemory_2_state_state <= _GEN_3551;
    end
    if (reset) begin
      TBEMemory_2_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'h2 == idxAlloc[3:0]) begin
        TBEMemory_2_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h2 == idxAlloc[3:0]) begin
          TBEMemory_2_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEMemory_2_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEMemory_2_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEMemory_2_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEMemory_2_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEMemory_2_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEMemory_2_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEMemory_2_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h2 == idxUpdate_0[3:0]) begin
                        TBEMemory_2_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEMemory_2_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEMemory_2_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h2 == idxUpdate_0[3:0]) begin
                        TBEMemory_2_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h2 == idxAlloc[3:0]) begin
                        TBEMemory_2_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'h2 == idxUpdate_0[3:0]) begin
                        TBEMemory_2_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h2 == idxUpdate_0[3:0]) begin
                          TBEMemory_2_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEMemory_2_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEMemory_2_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h2 == idxUpdate_0[3:0]) begin
                        TBEMemory_2_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_2_way <= _GEN_451;
                end
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEMemory_2_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_2_way <= _GEN_451;
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_way <= 3'h2;
                  end else begin
                    TBEMemory_2_way <= _GEN_451;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_2_way <= _GEN_451;
                  end else if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_2_way <= _GEN_451;
                  end
                end else begin
                  TBEMemory_2_way <= _GEN_451;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEMemory_2_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_2_way <= _GEN_451;
                    end
                  end else if (_T_111) begin
                    if (4'h2 == idxUpdate_1[3:0]) begin
                      TBEMemory_2_way <= 3'h2;
                    end else begin
                      TBEMemory_2_way <= _GEN_451;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_2_way <= _GEN_451;
                    end else if (4'h2 == idxUpdate_1[3:0]) begin
                      TBEMemory_2_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_2_way <= _GEN_451;
                    end
                  end else begin
                    TBEMemory_2_way <= _GEN_451;
                  end
                end else if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEMemory_2_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_2_way <= _GEN_451;
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_way <= 3'h2;
                  end else begin
                    TBEMemory_2_way <= _GEN_451;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_2_way <= _GEN_451;
                  end else if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_2_way <= _GEN_451;
                  end
                end else begin
                  TBEMemory_2_way <= _GEN_451;
                end
              end else begin
                TBEMemory_2_way <= _GEN_965;
              end
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEMemory_2_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_2_way <= _GEN_965;
                end
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_way <= 3'h2;
                end else begin
                  TBEMemory_2_way <= _GEN_965;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_2_way <= _GEN_965;
                end else if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_2_way <= _GEN_965;
                end
              end else begin
                TBEMemory_2_way <= _GEN_965;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEMemory_2_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_2_way <= _GEN_965;
                  end
                end else if (_T_133) begin
                  if (4'h2 == idxUpdate_2[3:0]) begin
                    TBEMemory_2_way <= 3'h2;
                  end else begin
                    TBEMemory_2_way <= _GEN_965;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_2_way <= _GEN_965;
                  end else if (4'h2 == idxUpdate_2[3:0]) begin
                    TBEMemory_2_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_2_way <= _GEN_965;
                  end
                end else begin
                  TBEMemory_2_way <= _GEN_965;
                end
              end else if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEMemory_2_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_2_way <= _GEN_965;
                end
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_way <= 3'h2;
                end else begin
                  TBEMemory_2_way <= _GEN_965;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_2_way <= _GEN_965;
                end else if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_2_way <= _GEN_965;
                end
              end else begin
                TBEMemory_2_way <= _GEN_965;
              end
            end else begin
              TBEMemory_2_way <= _GEN_1479;
            end
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEMemory_2_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_2_way <= _GEN_1479;
              end
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_way <= 3'h2;
              end else begin
                TBEMemory_2_way <= _GEN_1479;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_2_way <= _GEN_1479;
              end else if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_2_way <= _GEN_1479;
              end
            end else begin
              TBEMemory_2_way <= _GEN_1479;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEMemory_2_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_2_way <= _GEN_1479;
                end
              end else if (_T_155) begin
                if (4'h2 == idxUpdate_3[3:0]) begin
                  TBEMemory_2_way <= 3'h2;
                end else begin
                  TBEMemory_2_way <= _GEN_1479;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_2_way <= _GEN_1479;
                end else if (4'h2 == idxUpdate_3[3:0]) begin
                  TBEMemory_2_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_2_way <= _GEN_1479;
                end
              end else begin
                TBEMemory_2_way <= _GEN_1479;
              end
            end else if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEMemory_2_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_2_way <= _GEN_1479;
              end
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_way <= 3'h2;
              end else begin
                TBEMemory_2_way <= _GEN_1479;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_2_way <= _GEN_1479;
              end else if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_2_way <= _GEN_1479;
              end
            end else begin
              TBEMemory_2_way <= _GEN_1479;
            end
          end else begin
            TBEMemory_2_way <= _GEN_1993;
          end
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEMemory_2_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_2_way <= _GEN_1993;
            end
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_way <= 3'h2;
            end else begin
              TBEMemory_2_way <= _GEN_1993;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_2_way <= _GEN_1993;
            end else if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_2_way <= _GEN_1993;
            end
          end else begin
            TBEMemory_2_way <= _GEN_1993;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEMemory_2_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_2_way <= _GEN_1993;
              end
            end else if (_T_177) begin
              if (4'h2 == idxUpdate_4[3:0]) begin
                TBEMemory_2_way <= 3'h2;
              end else begin
                TBEMemory_2_way <= _GEN_1993;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_2_way <= _GEN_1993;
              end else if (4'h2 == idxUpdate_4[3:0]) begin
                TBEMemory_2_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_2_way <= _GEN_1993;
              end
            end else begin
              TBEMemory_2_way <= _GEN_1993;
            end
          end else if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEMemory_2_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_2_way <= _GEN_1993;
            end
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_way <= 3'h2;
            end else begin
              TBEMemory_2_way <= _GEN_1993;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_2_way <= _GEN_1993;
            end else if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_2_way <= _GEN_1993;
            end
          end else begin
            TBEMemory_2_way <= _GEN_1993;
          end
        end else begin
          TBEMemory_2_way <= _GEN_2507;
        end
      end else if (_T_221) begin
        if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEMemory_2_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_2_way <= _GEN_2507;
          end
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_way <= 3'h2;
          end else begin
            TBEMemory_2_way <= _GEN_2507;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_2_way <= _GEN_2507;
          end else if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_2_way <= _GEN_2507;
          end
        end else begin
          TBEMemory_2_way <= _GEN_2507;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEMemory_2_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_2_way <= _GEN_2507;
            end
          end else if (_T_199) begin
            if (4'h2 == idxUpdate_5[3:0]) begin
              TBEMemory_2_way <= 3'h2;
            end else begin
              TBEMemory_2_way <= _GEN_2507;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_2_way <= _GEN_2507;
            end else if (4'h2 == idxUpdate_5[3:0]) begin
              TBEMemory_2_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_2_way <= _GEN_2507;
            end
          end else begin
            TBEMemory_2_way <= _GEN_2507;
          end
        end else if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEMemory_2_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_2_way <= _GEN_2507;
          end
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_way <= 3'h2;
          end else begin
            TBEMemory_2_way <= _GEN_2507;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_2_way <= _GEN_2507;
          end else if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_2_way <= _GEN_2507;
          end
        end else begin
          TBEMemory_2_way <= _GEN_2507;
        end
      end else begin
        TBEMemory_2_way <= _GEN_3021;
      end
    end else if (_T_243) begin
      if (4'h2 == idxUpdate_7[3:0]) begin
        TBEMemory_2_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'h2 == idxAlloc[3:0]) begin
          TBEMemory_2_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_2_way <= _GEN_3021;
        end
      end else if (_T_221) begin
        if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_way <= 3'h2;
        end else begin
          TBEMemory_2_way <= _GEN_3021;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_2_way <= _GEN_3021;
        end else if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_2_way <= _GEN_3021;
        end
      end else begin
        TBEMemory_2_way <= _GEN_3021;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEMemory_2_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_2_way <= _GEN_3021;
          end
        end else if (_T_221) begin
          if (4'h2 == idxUpdate_6[3:0]) begin
            TBEMemory_2_way <= 3'h2;
          end else begin
            TBEMemory_2_way <= _GEN_3021;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_2_way <= _GEN_3021;
          end else if (4'h2 == idxUpdate_6[3:0]) begin
            TBEMemory_2_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_2_way <= _GEN_3021;
          end
        end else begin
          TBEMemory_2_way <= _GEN_3021;
        end
      end else if (4'h2 == idxUpdate_7[3:0]) begin
        TBEMemory_2_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h2 == idxAlloc[3:0]) begin
          TBEMemory_2_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_2_way <= _GEN_3021;
        end
      end else if (_T_221) begin
        if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_way <= 3'h2;
        end else begin
          TBEMemory_2_way <= _GEN_3021;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_2_way <= _GEN_3021;
        end else if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_2_way <= _GEN_3021;
        end
      end else begin
        TBEMemory_2_way <= _GEN_3021;
      end
    end else begin
      TBEMemory_2_way <= _GEN_3535;
    end
    if (reset) begin
      TBEMemory_2_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h2 == idxAlloc[3:0]) begin
        TBEMemory_2_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'h2 == idxAlloc[3:0]) begin
          TBEMemory_2_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEMemory_2_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEMemory_2_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEMemory_2_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEMemory_2_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEMemory_2_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEMemory_2_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEMemory_2_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h2 == idxUpdate_0[3:0]) begin
                        TBEMemory_2_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEMemory_2_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEMemory_2_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h2 == idxUpdate_0[3:0]) begin
                        TBEMemory_2_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h2 == idxUpdate_1[3:0]) begin
                      TBEMemory_2_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'h2 == idxAlloc[3:0]) begin
                        TBEMemory_2_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'h2 == idxUpdate_0[3:0]) begin
                        TBEMemory_2_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'h2 == idxUpdate_0[3:0]) begin
                          TBEMemory_2_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEMemory_2_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEMemory_2_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h2 == idxUpdate_0[3:0]) begin
                        TBEMemory_2_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_435;
                end
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEMemory_2_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_435;
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_435;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h2 == idxUpdate_1[3:0]) begin
                      TBEMemory_2_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_2_fields_0 <= _GEN_435;
                    end
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_435;
                  end
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_435;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h2 == idxUpdate_2[3:0]) begin
                    TBEMemory_2_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEMemory_2_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_2_fields_0 <= _GEN_435;
                    end
                  end else if (_T_111) begin
                    if (4'h2 == idxUpdate_1[3:0]) begin
                      TBEMemory_2_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_2_fields_0 <= _GEN_435;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'h2 == idxUpdate_1[3:0]) begin
                        TBEMemory_2_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_2_fields_0 <= _GEN_435;
                      end
                    end else begin
                      TBEMemory_2_fields_0 <= _GEN_435;
                    end
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_435;
                  end
                end else if (isAlloc_1) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEMemory_2_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_435;
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEMemory_2_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_435;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h2 == idxUpdate_1[3:0]) begin
                      TBEMemory_2_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_2_fields_0 <= _GEN_435;
                    end
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_435;
                  end
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_435;
                end
              end else begin
                TBEMemory_2_fields_0 <= _GEN_949;
              end
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEMemory_2_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_949;
                end
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_949;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h2 == idxUpdate_2[3:0]) begin
                    TBEMemory_2_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_949;
                  end
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_949;
                end
              end else begin
                TBEMemory_2_fields_0 <= _GEN_949;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h2 == idxUpdate_3[3:0]) begin
                  TBEMemory_2_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEMemory_2_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_949;
                  end
                end else if (_T_133) begin
                  if (4'h2 == idxUpdate_2[3:0]) begin
                    TBEMemory_2_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_949;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'h2 == idxUpdate_2[3:0]) begin
                      TBEMemory_2_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_2_fields_0 <= _GEN_949;
                    end
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_949;
                  end
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_949;
                end
              end else if (isAlloc_2) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEMemory_2_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_949;
                end
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEMemory_2_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_949;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h2 == idxUpdate_2[3:0]) begin
                    TBEMemory_2_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_949;
                  end
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_949;
                end
              end else begin
                TBEMemory_2_fields_0 <= _GEN_949;
              end
            end else begin
              TBEMemory_2_fields_0 <= _GEN_1463;
            end
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEMemory_2_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_2_fields_0 <= _GEN_1463;
              end
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_fields_0 <= 32'h0;
              end else begin
                TBEMemory_2_fields_0 <= _GEN_1463;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h2 == idxUpdate_3[3:0]) begin
                  TBEMemory_2_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_1463;
                end
              end else begin
                TBEMemory_2_fields_0 <= _GEN_1463;
              end
            end else begin
              TBEMemory_2_fields_0 <= _GEN_1463;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h2 == idxUpdate_4[3:0]) begin
                TBEMemory_2_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEMemory_2_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_1463;
                end
              end else if (_T_155) begin
                if (4'h2 == idxUpdate_3[3:0]) begin
                  TBEMemory_2_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_1463;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'h2 == idxUpdate_3[3:0]) begin
                    TBEMemory_2_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_2_fields_0 <= _GEN_1463;
                  end
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_1463;
                end
              end else begin
                TBEMemory_2_fields_0 <= _GEN_1463;
              end
            end else if (isAlloc_3) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEMemory_2_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_2_fields_0 <= _GEN_1463;
              end
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEMemory_2_fields_0 <= 32'h0;
              end else begin
                TBEMemory_2_fields_0 <= _GEN_1463;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h2 == idxUpdate_3[3:0]) begin
                  TBEMemory_2_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_1463;
                end
              end else begin
                TBEMemory_2_fields_0 <= _GEN_1463;
              end
            end else begin
              TBEMemory_2_fields_0 <= _GEN_1463;
            end
          end else begin
            TBEMemory_2_fields_0 <= _GEN_1977;
          end
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEMemory_2_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_2_fields_0 <= _GEN_1977;
            end
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_fields_0 <= 32'h0;
            end else begin
              TBEMemory_2_fields_0 <= _GEN_1977;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h2 == idxUpdate_4[3:0]) begin
                TBEMemory_2_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_2_fields_0 <= _GEN_1977;
              end
            end else begin
              TBEMemory_2_fields_0 <= _GEN_1977;
            end
          end else begin
            TBEMemory_2_fields_0 <= _GEN_1977;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h2 == idxUpdate_5[3:0]) begin
              TBEMemory_2_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEMemory_2_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_2_fields_0 <= _GEN_1977;
              end
            end else if (_T_177) begin
              if (4'h2 == idxUpdate_4[3:0]) begin
                TBEMemory_2_fields_0 <= 32'h0;
              end else begin
                TBEMemory_2_fields_0 <= _GEN_1977;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'h2 == idxUpdate_4[3:0]) begin
                  TBEMemory_2_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_2_fields_0 <= _GEN_1977;
                end
              end else begin
                TBEMemory_2_fields_0 <= _GEN_1977;
              end
            end else begin
              TBEMemory_2_fields_0 <= _GEN_1977;
            end
          end else if (isAlloc_4) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEMemory_2_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_2_fields_0 <= _GEN_1977;
            end
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEMemory_2_fields_0 <= 32'h0;
            end else begin
              TBEMemory_2_fields_0 <= _GEN_1977;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h2 == idxUpdate_4[3:0]) begin
                TBEMemory_2_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_2_fields_0 <= _GEN_1977;
              end
            end else begin
              TBEMemory_2_fields_0 <= _GEN_1977;
            end
          end else begin
            TBEMemory_2_fields_0 <= _GEN_1977;
          end
        end else begin
          TBEMemory_2_fields_0 <= _GEN_2491;
        end
      end else if (_T_221) begin
        if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEMemory_2_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_2_fields_0 <= _GEN_2491;
          end
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_fields_0 <= 32'h0;
          end else begin
            TBEMemory_2_fields_0 <= _GEN_2491;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h2 == idxUpdate_5[3:0]) begin
              TBEMemory_2_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_2_fields_0 <= _GEN_2491;
            end
          end else begin
            TBEMemory_2_fields_0 <= _GEN_2491;
          end
        end else begin
          TBEMemory_2_fields_0 <= _GEN_2491;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h2 == idxUpdate_6[3:0]) begin
            TBEMemory_2_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEMemory_2_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_2_fields_0 <= _GEN_2491;
            end
          end else if (_T_199) begin
            if (4'h2 == idxUpdate_5[3:0]) begin
              TBEMemory_2_fields_0 <= 32'h0;
            end else begin
              TBEMemory_2_fields_0 <= _GEN_2491;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'h2 == idxUpdate_5[3:0]) begin
                TBEMemory_2_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_2_fields_0 <= _GEN_2491;
              end
            end else begin
              TBEMemory_2_fields_0 <= _GEN_2491;
            end
          end else begin
            TBEMemory_2_fields_0 <= _GEN_2491;
          end
        end else if (isAlloc_5) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEMemory_2_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_2_fields_0 <= _GEN_2491;
          end
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEMemory_2_fields_0 <= 32'h0;
          end else begin
            TBEMemory_2_fields_0 <= _GEN_2491;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h2 == idxUpdate_5[3:0]) begin
              TBEMemory_2_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_2_fields_0 <= _GEN_2491;
            end
          end else begin
            TBEMemory_2_fields_0 <= _GEN_2491;
          end
        end else begin
          TBEMemory_2_fields_0 <= _GEN_2491;
        end
      end else begin
        TBEMemory_2_fields_0 <= _GEN_3005;
      end
    end else if (_T_243) begin
      if (4'h2 == idxUpdate_7[3:0]) begin
        TBEMemory_2_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h2 == idxAlloc[3:0]) begin
          TBEMemory_2_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_2_fields_0 <= _GEN_3005;
        end
      end else if (_T_221) begin
        if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_fields_0 <= 32'h0;
        end else begin
          TBEMemory_2_fields_0 <= _GEN_3005;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h2 == idxUpdate_6[3:0]) begin
            TBEMemory_2_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_2_fields_0 <= _GEN_3005;
          end
        end else begin
          TBEMemory_2_fields_0 <= _GEN_3005;
        end
      end else begin
        TBEMemory_2_fields_0 <= _GEN_3005;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'h2 == idxUpdate_7[3:0]) begin
          TBEMemory_2_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEMemory_2_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_2_fields_0 <= _GEN_3005;
          end
        end else if (_T_221) begin
          if (4'h2 == idxUpdate_6[3:0]) begin
            TBEMemory_2_fields_0 <= 32'h0;
          end else begin
            TBEMemory_2_fields_0 <= _GEN_3005;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'h2 == idxUpdate_6[3:0]) begin
              TBEMemory_2_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_2_fields_0 <= _GEN_3005;
            end
          end else begin
            TBEMemory_2_fields_0 <= _GEN_3005;
          end
        end else begin
          TBEMemory_2_fields_0 <= _GEN_3005;
        end
      end else if (isAlloc_6) begin
        if (4'h2 == idxAlloc[3:0]) begin
          TBEMemory_2_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_2_fields_0 <= _GEN_3005;
        end
      end else if (_T_221) begin
        if (4'h2 == idxUpdate_6[3:0]) begin
          TBEMemory_2_fields_0 <= 32'h0;
        end else begin
          TBEMemory_2_fields_0 <= _GEN_3005;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h2 == idxUpdate_6[3:0]) begin
            TBEMemory_2_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_2_fields_0 <= _GEN_3005;
          end
        end else begin
          TBEMemory_2_fields_0 <= _GEN_3005;
        end
      end else begin
        TBEMemory_2_fields_0 <= _GEN_3005;
      end
    end else begin
      TBEMemory_2_fields_0 <= _GEN_3519;
    end
    if (reset) begin
      TBEMemory_3_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'h3 == idxAlloc[3:0]) begin
        TBEMemory_3_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h3 == idxAlloc[3:0]) begin
          TBEMemory_3_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEMemory_3_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEMemory_3_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEMemory_3_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEMemory_3_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEMemory_3_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEMemory_3_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEMemory_3_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h3 == idxUpdate_0[3:0]) begin
                        TBEMemory_3_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEMemory_3_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEMemory_3_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h3 == idxUpdate_0[3:0]) begin
                        TBEMemory_3_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h3 == idxAlloc[3:0]) begin
                        TBEMemory_3_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'h3 == idxUpdate_0[3:0]) begin
                        TBEMemory_3_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h3 == idxUpdate_0[3:0]) begin
                          TBEMemory_3_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEMemory_3_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEMemory_3_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h3 == idxUpdate_0[3:0]) begin
                        TBEMemory_3_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_3_state_state <= _GEN_468;
                end
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEMemory_3_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_3_state_state <= _GEN_468;
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_state_state <= 2'h0;
                  end else begin
                    TBEMemory_3_state_state <= _GEN_468;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_3_state_state <= _GEN_468;
                  end else if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_3_state_state <= _GEN_468;
                  end
                end else begin
                  TBEMemory_3_state_state <= _GEN_468;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEMemory_3_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_3_state_state <= _GEN_468;
                    end
                  end else if (_T_111) begin
                    if (4'h3 == idxUpdate_1[3:0]) begin
                      TBEMemory_3_state_state <= 2'h0;
                    end else begin
                      TBEMemory_3_state_state <= _GEN_468;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_3_state_state <= _GEN_468;
                    end else if (4'h3 == idxUpdate_1[3:0]) begin
                      TBEMemory_3_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_3_state_state <= _GEN_468;
                    end
                  end else begin
                    TBEMemory_3_state_state <= _GEN_468;
                  end
                end else if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEMemory_3_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_3_state_state <= _GEN_468;
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_state_state <= 2'h0;
                  end else begin
                    TBEMemory_3_state_state <= _GEN_468;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_3_state_state <= _GEN_468;
                  end else if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_3_state_state <= _GEN_468;
                  end
                end else begin
                  TBEMemory_3_state_state <= _GEN_468;
                end
              end else begin
                TBEMemory_3_state_state <= _GEN_982;
              end
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEMemory_3_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_3_state_state <= _GEN_982;
                end
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_state_state <= 2'h0;
                end else begin
                  TBEMemory_3_state_state <= _GEN_982;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_3_state_state <= _GEN_982;
                end else if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_3_state_state <= _GEN_982;
                end
              end else begin
                TBEMemory_3_state_state <= _GEN_982;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEMemory_3_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_3_state_state <= _GEN_982;
                  end
                end else if (_T_133) begin
                  if (4'h3 == idxUpdate_2[3:0]) begin
                    TBEMemory_3_state_state <= 2'h0;
                  end else begin
                    TBEMemory_3_state_state <= _GEN_982;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_3_state_state <= _GEN_982;
                  end else if (4'h3 == idxUpdate_2[3:0]) begin
                    TBEMemory_3_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_3_state_state <= _GEN_982;
                  end
                end else begin
                  TBEMemory_3_state_state <= _GEN_982;
                end
              end else if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEMemory_3_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_3_state_state <= _GEN_982;
                end
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_state_state <= 2'h0;
                end else begin
                  TBEMemory_3_state_state <= _GEN_982;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_3_state_state <= _GEN_982;
                end else if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_3_state_state <= _GEN_982;
                end
              end else begin
                TBEMemory_3_state_state <= _GEN_982;
              end
            end else begin
              TBEMemory_3_state_state <= _GEN_1496;
            end
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEMemory_3_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_3_state_state <= _GEN_1496;
              end
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_state_state <= 2'h0;
              end else begin
                TBEMemory_3_state_state <= _GEN_1496;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_3_state_state <= _GEN_1496;
              end else if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_3_state_state <= _GEN_1496;
              end
            end else begin
              TBEMemory_3_state_state <= _GEN_1496;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEMemory_3_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_3_state_state <= _GEN_1496;
                end
              end else if (_T_155) begin
                if (4'h3 == idxUpdate_3[3:0]) begin
                  TBEMemory_3_state_state <= 2'h0;
                end else begin
                  TBEMemory_3_state_state <= _GEN_1496;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_3_state_state <= _GEN_1496;
                end else if (4'h3 == idxUpdate_3[3:0]) begin
                  TBEMemory_3_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_3_state_state <= _GEN_1496;
                end
              end else begin
                TBEMemory_3_state_state <= _GEN_1496;
              end
            end else if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEMemory_3_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_3_state_state <= _GEN_1496;
              end
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_state_state <= 2'h0;
              end else begin
                TBEMemory_3_state_state <= _GEN_1496;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_3_state_state <= _GEN_1496;
              end else if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_3_state_state <= _GEN_1496;
              end
            end else begin
              TBEMemory_3_state_state <= _GEN_1496;
            end
          end else begin
            TBEMemory_3_state_state <= _GEN_2010;
          end
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEMemory_3_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_3_state_state <= _GEN_2010;
            end
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_state_state <= 2'h0;
            end else begin
              TBEMemory_3_state_state <= _GEN_2010;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_3_state_state <= _GEN_2010;
            end else if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_3_state_state <= _GEN_2010;
            end
          end else begin
            TBEMemory_3_state_state <= _GEN_2010;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEMemory_3_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_3_state_state <= _GEN_2010;
              end
            end else if (_T_177) begin
              if (4'h3 == idxUpdate_4[3:0]) begin
                TBEMemory_3_state_state <= 2'h0;
              end else begin
                TBEMemory_3_state_state <= _GEN_2010;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_3_state_state <= _GEN_2010;
              end else if (4'h3 == idxUpdate_4[3:0]) begin
                TBEMemory_3_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_3_state_state <= _GEN_2010;
              end
            end else begin
              TBEMemory_3_state_state <= _GEN_2010;
            end
          end else if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEMemory_3_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_3_state_state <= _GEN_2010;
            end
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_state_state <= 2'h0;
            end else begin
              TBEMemory_3_state_state <= _GEN_2010;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_3_state_state <= _GEN_2010;
            end else if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_3_state_state <= _GEN_2010;
            end
          end else begin
            TBEMemory_3_state_state <= _GEN_2010;
          end
        end else begin
          TBEMemory_3_state_state <= _GEN_2524;
        end
      end else if (_T_221) begin
        if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEMemory_3_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_3_state_state <= _GEN_2524;
          end
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_state_state <= 2'h0;
          end else begin
            TBEMemory_3_state_state <= _GEN_2524;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_3_state_state <= _GEN_2524;
          end else if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_3_state_state <= _GEN_2524;
          end
        end else begin
          TBEMemory_3_state_state <= _GEN_2524;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEMemory_3_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_3_state_state <= _GEN_2524;
            end
          end else if (_T_199) begin
            if (4'h3 == idxUpdate_5[3:0]) begin
              TBEMemory_3_state_state <= 2'h0;
            end else begin
              TBEMemory_3_state_state <= _GEN_2524;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_3_state_state <= _GEN_2524;
            end else if (4'h3 == idxUpdate_5[3:0]) begin
              TBEMemory_3_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_3_state_state <= _GEN_2524;
            end
          end else begin
            TBEMemory_3_state_state <= _GEN_2524;
          end
        end else if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEMemory_3_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_3_state_state <= _GEN_2524;
          end
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_state_state <= 2'h0;
          end else begin
            TBEMemory_3_state_state <= _GEN_2524;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_3_state_state <= _GEN_2524;
          end else if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_3_state_state <= _GEN_2524;
          end
        end else begin
          TBEMemory_3_state_state <= _GEN_2524;
        end
      end else begin
        TBEMemory_3_state_state <= _GEN_3038;
      end
    end else if (_T_243) begin
      if (4'h3 == idxUpdate_7[3:0]) begin
        TBEMemory_3_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'h3 == idxAlloc[3:0]) begin
          TBEMemory_3_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_3_state_state <= _GEN_3038;
        end
      end else if (_T_221) begin
        if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_state_state <= 2'h0;
        end else begin
          TBEMemory_3_state_state <= _GEN_3038;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_3_state_state <= _GEN_3038;
        end else if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_3_state_state <= _GEN_3038;
        end
      end else begin
        TBEMemory_3_state_state <= _GEN_3038;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEMemory_3_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_3_state_state <= _GEN_3038;
          end
        end else if (_T_221) begin
          if (4'h3 == idxUpdate_6[3:0]) begin
            TBEMemory_3_state_state <= 2'h0;
          end else begin
            TBEMemory_3_state_state <= _GEN_3038;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_3_state_state <= _GEN_3038;
          end else if (4'h3 == idxUpdate_6[3:0]) begin
            TBEMemory_3_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_3_state_state <= _GEN_3038;
          end
        end else begin
          TBEMemory_3_state_state <= _GEN_3038;
        end
      end else if (4'h3 == idxUpdate_7[3:0]) begin
        TBEMemory_3_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h3 == idxAlloc[3:0]) begin
          TBEMemory_3_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_3_state_state <= _GEN_3038;
        end
      end else if (_T_221) begin
        if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_state_state <= 2'h0;
        end else begin
          TBEMemory_3_state_state <= _GEN_3038;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_3_state_state <= _GEN_3038;
        end else if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_3_state_state <= _GEN_3038;
        end
      end else begin
        TBEMemory_3_state_state <= _GEN_3038;
      end
    end else begin
      TBEMemory_3_state_state <= _GEN_3552;
    end
    if (reset) begin
      TBEMemory_3_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'h3 == idxAlloc[3:0]) begin
        TBEMemory_3_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h3 == idxAlloc[3:0]) begin
          TBEMemory_3_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEMemory_3_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEMemory_3_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEMemory_3_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEMemory_3_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEMemory_3_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEMemory_3_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEMemory_3_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h3 == idxUpdate_0[3:0]) begin
                        TBEMemory_3_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEMemory_3_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEMemory_3_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h3 == idxUpdate_0[3:0]) begin
                        TBEMemory_3_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h3 == idxAlloc[3:0]) begin
                        TBEMemory_3_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'h3 == idxUpdate_0[3:0]) begin
                        TBEMemory_3_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h3 == idxUpdate_0[3:0]) begin
                          TBEMemory_3_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEMemory_3_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEMemory_3_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h3 == idxUpdate_0[3:0]) begin
                        TBEMemory_3_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_3_way <= _GEN_452;
                end
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEMemory_3_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_3_way <= _GEN_452;
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_way <= 3'h2;
                  end else begin
                    TBEMemory_3_way <= _GEN_452;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_3_way <= _GEN_452;
                  end else if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_3_way <= _GEN_452;
                  end
                end else begin
                  TBEMemory_3_way <= _GEN_452;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEMemory_3_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_3_way <= _GEN_452;
                    end
                  end else if (_T_111) begin
                    if (4'h3 == idxUpdate_1[3:0]) begin
                      TBEMemory_3_way <= 3'h2;
                    end else begin
                      TBEMemory_3_way <= _GEN_452;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_3_way <= _GEN_452;
                    end else if (4'h3 == idxUpdate_1[3:0]) begin
                      TBEMemory_3_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_3_way <= _GEN_452;
                    end
                  end else begin
                    TBEMemory_3_way <= _GEN_452;
                  end
                end else if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEMemory_3_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_3_way <= _GEN_452;
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_way <= 3'h2;
                  end else begin
                    TBEMemory_3_way <= _GEN_452;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_3_way <= _GEN_452;
                  end else if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_3_way <= _GEN_452;
                  end
                end else begin
                  TBEMemory_3_way <= _GEN_452;
                end
              end else begin
                TBEMemory_3_way <= _GEN_966;
              end
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEMemory_3_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_3_way <= _GEN_966;
                end
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_way <= 3'h2;
                end else begin
                  TBEMemory_3_way <= _GEN_966;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_3_way <= _GEN_966;
                end else if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_3_way <= _GEN_966;
                end
              end else begin
                TBEMemory_3_way <= _GEN_966;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEMemory_3_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_3_way <= _GEN_966;
                  end
                end else if (_T_133) begin
                  if (4'h3 == idxUpdate_2[3:0]) begin
                    TBEMemory_3_way <= 3'h2;
                  end else begin
                    TBEMemory_3_way <= _GEN_966;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_3_way <= _GEN_966;
                  end else if (4'h3 == idxUpdate_2[3:0]) begin
                    TBEMemory_3_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_3_way <= _GEN_966;
                  end
                end else begin
                  TBEMemory_3_way <= _GEN_966;
                end
              end else if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEMemory_3_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_3_way <= _GEN_966;
                end
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_way <= 3'h2;
                end else begin
                  TBEMemory_3_way <= _GEN_966;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_3_way <= _GEN_966;
                end else if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_3_way <= _GEN_966;
                end
              end else begin
                TBEMemory_3_way <= _GEN_966;
              end
            end else begin
              TBEMemory_3_way <= _GEN_1480;
            end
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEMemory_3_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_3_way <= _GEN_1480;
              end
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_way <= 3'h2;
              end else begin
                TBEMemory_3_way <= _GEN_1480;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_3_way <= _GEN_1480;
              end else if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_3_way <= _GEN_1480;
              end
            end else begin
              TBEMemory_3_way <= _GEN_1480;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEMemory_3_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_3_way <= _GEN_1480;
                end
              end else if (_T_155) begin
                if (4'h3 == idxUpdate_3[3:0]) begin
                  TBEMemory_3_way <= 3'h2;
                end else begin
                  TBEMemory_3_way <= _GEN_1480;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_3_way <= _GEN_1480;
                end else if (4'h3 == idxUpdate_3[3:0]) begin
                  TBEMemory_3_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_3_way <= _GEN_1480;
                end
              end else begin
                TBEMemory_3_way <= _GEN_1480;
              end
            end else if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEMemory_3_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_3_way <= _GEN_1480;
              end
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_way <= 3'h2;
              end else begin
                TBEMemory_3_way <= _GEN_1480;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_3_way <= _GEN_1480;
              end else if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_3_way <= _GEN_1480;
              end
            end else begin
              TBEMemory_3_way <= _GEN_1480;
            end
          end else begin
            TBEMemory_3_way <= _GEN_1994;
          end
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEMemory_3_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_3_way <= _GEN_1994;
            end
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_way <= 3'h2;
            end else begin
              TBEMemory_3_way <= _GEN_1994;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_3_way <= _GEN_1994;
            end else if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_3_way <= _GEN_1994;
            end
          end else begin
            TBEMemory_3_way <= _GEN_1994;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEMemory_3_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_3_way <= _GEN_1994;
              end
            end else if (_T_177) begin
              if (4'h3 == idxUpdate_4[3:0]) begin
                TBEMemory_3_way <= 3'h2;
              end else begin
                TBEMemory_3_way <= _GEN_1994;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_3_way <= _GEN_1994;
              end else if (4'h3 == idxUpdate_4[3:0]) begin
                TBEMemory_3_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_3_way <= _GEN_1994;
              end
            end else begin
              TBEMemory_3_way <= _GEN_1994;
            end
          end else if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEMemory_3_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_3_way <= _GEN_1994;
            end
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_way <= 3'h2;
            end else begin
              TBEMemory_3_way <= _GEN_1994;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_3_way <= _GEN_1994;
            end else if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_3_way <= _GEN_1994;
            end
          end else begin
            TBEMemory_3_way <= _GEN_1994;
          end
        end else begin
          TBEMemory_3_way <= _GEN_2508;
        end
      end else if (_T_221) begin
        if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEMemory_3_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_3_way <= _GEN_2508;
          end
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_way <= 3'h2;
          end else begin
            TBEMemory_3_way <= _GEN_2508;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_3_way <= _GEN_2508;
          end else if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_3_way <= _GEN_2508;
          end
        end else begin
          TBEMemory_3_way <= _GEN_2508;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEMemory_3_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_3_way <= _GEN_2508;
            end
          end else if (_T_199) begin
            if (4'h3 == idxUpdate_5[3:0]) begin
              TBEMemory_3_way <= 3'h2;
            end else begin
              TBEMemory_3_way <= _GEN_2508;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_3_way <= _GEN_2508;
            end else if (4'h3 == idxUpdate_5[3:0]) begin
              TBEMemory_3_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_3_way <= _GEN_2508;
            end
          end else begin
            TBEMemory_3_way <= _GEN_2508;
          end
        end else if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEMemory_3_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_3_way <= _GEN_2508;
          end
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_way <= 3'h2;
          end else begin
            TBEMemory_3_way <= _GEN_2508;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_3_way <= _GEN_2508;
          end else if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_3_way <= _GEN_2508;
          end
        end else begin
          TBEMemory_3_way <= _GEN_2508;
        end
      end else begin
        TBEMemory_3_way <= _GEN_3022;
      end
    end else if (_T_243) begin
      if (4'h3 == idxUpdate_7[3:0]) begin
        TBEMemory_3_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'h3 == idxAlloc[3:0]) begin
          TBEMemory_3_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_3_way <= _GEN_3022;
        end
      end else if (_T_221) begin
        if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_way <= 3'h2;
        end else begin
          TBEMemory_3_way <= _GEN_3022;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_3_way <= _GEN_3022;
        end else if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_3_way <= _GEN_3022;
        end
      end else begin
        TBEMemory_3_way <= _GEN_3022;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEMemory_3_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_3_way <= _GEN_3022;
          end
        end else if (_T_221) begin
          if (4'h3 == idxUpdate_6[3:0]) begin
            TBEMemory_3_way <= 3'h2;
          end else begin
            TBEMemory_3_way <= _GEN_3022;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_3_way <= _GEN_3022;
          end else if (4'h3 == idxUpdate_6[3:0]) begin
            TBEMemory_3_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_3_way <= _GEN_3022;
          end
        end else begin
          TBEMemory_3_way <= _GEN_3022;
        end
      end else if (4'h3 == idxUpdate_7[3:0]) begin
        TBEMemory_3_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h3 == idxAlloc[3:0]) begin
          TBEMemory_3_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_3_way <= _GEN_3022;
        end
      end else if (_T_221) begin
        if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_way <= 3'h2;
        end else begin
          TBEMemory_3_way <= _GEN_3022;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_3_way <= _GEN_3022;
        end else if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_3_way <= _GEN_3022;
        end
      end else begin
        TBEMemory_3_way <= _GEN_3022;
      end
    end else begin
      TBEMemory_3_way <= _GEN_3536;
    end
    if (reset) begin
      TBEMemory_3_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h3 == idxAlloc[3:0]) begin
        TBEMemory_3_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'h3 == idxAlloc[3:0]) begin
          TBEMemory_3_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEMemory_3_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEMemory_3_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEMemory_3_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEMemory_3_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEMemory_3_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEMemory_3_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEMemory_3_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h3 == idxUpdate_0[3:0]) begin
                        TBEMemory_3_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEMemory_3_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEMemory_3_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h3 == idxUpdate_0[3:0]) begin
                        TBEMemory_3_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h3 == idxUpdate_1[3:0]) begin
                      TBEMemory_3_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'h3 == idxAlloc[3:0]) begin
                        TBEMemory_3_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'h3 == idxUpdate_0[3:0]) begin
                        TBEMemory_3_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'h3 == idxUpdate_0[3:0]) begin
                          TBEMemory_3_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEMemory_3_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEMemory_3_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h3 == idxUpdate_0[3:0]) begin
                        TBEMemory_3_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_436;
                end
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEMemory_3_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_436;
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_436;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h3 == idxUpdate_1[3:0]) begin
                      TBEMemory_3_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_3_fields_0 <= _GEN_436;
                    end
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_436;
                  end
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_436;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h3 == idxUpdate_2[3:0]) begin
                    TBEMemory_3_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEMemory_3_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_3_fields_0 <= _GEN_436;
                    end
                  end else if (_T_111) begin
                    if (4'h3 == idxUpdate_1[3:0]) begin
                      TBEMemory_3_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_3_fields_0 <= _GEN_436;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'h3 == idxUpdate_1[3:0]) begin
                        TBEMemory_3_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_3_fields_0 <= _GEN_436;
                      end
                    end else begin
                      TBEMemory_3_fields_0 <= _GEN_436;
                    end
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_436;
                  end
                end else if (isAlloc_1) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEMemory_3_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_436;
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEMemory_3_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_436;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h3 == idxUpdate_1[3:0]) begin
                      TBEMemory_3_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_3_fields_0 <= _GEN_436;
                    end
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_436;
                  end
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_436;
                end
              end else begin
                TBEMemory_3_fields_0 <= _GEN_950;
              end
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEMemory_3_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_950;
                end
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_950;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h3 == idxUpdate_2[3:0]) begin
                    TBEMemory_3_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_950;
                  end
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_950;
                end
              end else begin
                TBEMemory_3_fields_0 <= _GEN_950;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h3 == idxUpdate_3[3:0]) begin
                  TBEMemory_3_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEMemory_3_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_950;
                  end
                end else if (_T_133) begin
                  if (4'h3 == idxUpdate_2[3:0]) begin
                    TBEMemory_3_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_950;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'h3 == idxUpdate_2[3:0]) begin
                      TBEMemory_3_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_3_fields_0 <= _GEN_950;
                    end
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_950;
                  end
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_950;
                end
              end else if (isAlloc_2) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEMemory_3_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_950;
                end
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEMemory_3_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_950;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h3 == idxUpdate_2[3:0]) begin
                    TBEMemory_3_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_950;
                  end
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_950;
                end
              end else begin
                TBEMemory_3_fields_0 <= _GEN_950;
              end
            end else begin
              TBEMemory_3_fields_0 <= _GEN_1464;
            end
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEMemory_3_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_3_fields_0 <= _GEN_1464;
              end
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_fields_0 <= 32'h0;
              end else begin
                TBEMemory_3_fields_0 <= _GEN_1464;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h3 == idxUpdate_3[3:0]) begin
                  TBEMemory_3_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_1464;
                end
              end else begin
                TBEMemory_3_fields_0 <= _GEN_1464;
              end
            end else begin
              TBEMemory_3_fields_0 <= _GEN_1464;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h3 == idxUpdate_4[3:0]) begin
                TBEMemory_3_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEMemory_3_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_1464;
                end
              end else if (_T_155) begin
                if (4'h3 == idxUpdate_3[3:0]) begin
                  TBEMemory_3_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_1464;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'h3 == idxUpdate_3[3:0]) begin
                    TBEMemory_3_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_3_fields_0 <= _GEN_1464;
                  end
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_1464;
                end
              end else begin
                TBEMemory_3_fields_0 <= _GEN_1464;
              end
            end else if (isAlloc_3) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEMemory_3_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_3_fields_0 <= _GEN_1464;
              end
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEMemory_3_fields_0 <= 32'h0;
              end else begin
                TBEMemory_3_fields_0 <= _GEN_1464;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h3 == idxUpdate_3[3:0]) begin
                  TBEMemory_3_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_1464;
                end
              end else begin
                TBEMemory_3_fields_0 <= _GEN_1464;
              end
            end else begin
              TBEMemory_3_fields_0 <= _GEN_1464;
            end
          end else begin
            TBEMemory_3_fields_0 <= _GEN_1978;
          end
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEMemory_3_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_3_fields_0 <= _GEN_1978;
            end
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_fields_0 <= 32'h0;
            end else begin
              TBEMemory_3_fields_0 <= _GEN_1978;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h3 == idxUpdate_4[3:0]) begin
                TBEMemory_3_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_3_fields_0 <= _GEN_1978;
              end
            end else begin
              TBEMemory_3_fields_0 <= _GEN_1978;
            end
          end else begin
            TBEMemory_3_fields_0 <= _GEN_1978;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h3 == idxUpdate_5[3:0]) begin
              TBEMemory_3_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEMemory_3_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_3_fields_0 <= _GEN_1978;
              end
            end else if (_T_177) begin
              if (4'h3 == idxUpdate_4[3:0]) begin
                TBEMemory_3_fields_0 <= 32'h0;
              end else begin
                TBEMemory_3_fields_0 <= _GEN_1978;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'h3 == idxUpdate_4[3:0]) begin
                  TBEMemory_3_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_3_fields_0 <= _GEN_1978;
                end
              end else begin
                TBEMemory_3_fields_0 <= _GEN_1978;
              end
            end else begin
              TBEMemory_3_fields_0 <= _GEN_1978;
            end
          end else if (isAlloc_4) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEMemory_3_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_3_fields_0 <= _GEN_1978;
            end
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEMemory_3_fields_0 <= 32'h0;
            end else begin
              TBEMemory_3_fields_0 <= _GEN_1978;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h3 == idxUpdate_4[3:0]) begin
                TBEMemory_3_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_3_fields_0 <= _GEN_1978;
              end
            end else begin
              TBEMemory_3_fields_0 <= _GEN_1978;
            end
          end else begin
            TBEMemory_3_fields_0 <= _GEN_1978;
          end
        end else begin
          TBEMemory_3_fields_0 <= _GEN_2492;
        end
      end else if (_T_221) begin
        if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEMemory_3_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_3_fields_0 <= _GEN_2492;
          end
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_fields_0 <= 32'h0;
          end else begin
            TBEMemory_3_fields_0 <= _GEN_2492;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h3 == idxUpdate_5[3:0]) begin
              TBEMemory_3_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_3_fields_0 <= _GEN_2492;
            end
          end else begin
            TBEMemory_3_fields_0 <= _GEN_2492;
          end
        end else begin
          TBEMemory_3_fields_0 <= _GEN_2492;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h3 == idxUpdate_6[3:0]) begin
            TBEMemory_3_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEMemory_3_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_3_fields_0 <= _GEN_2492;
            end
          end else if (_T_199) begin
            if (4'h3 == idxUpdate_5[3:0]) begin
              TBEMemory_3_fields_0 <= 32'h0;
            end else begin
              TBEMemory_3_fields_0 <= _GEN_2492;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'h3 == idxUpdate_5[3:0]) begin
                TBEMemory_3_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_3_fields_0 <= _GEN_2492;
              end
            end else begin
              TBEMemory_3_fields_0 <= _GEN_2492;
            end
          end else begin
            TBEMemory_3_fields_0 <= _GEN_2492;
          end
        end else if (isAlloc_5) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEMemory_3_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_3_fields_0 <= _GEN_2492;
          end
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEMemory_3_fields_0 <= 32'h0;
          end else begin
            TBEMemory_3_fields_0 <= _GEN_2492;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h3 == idxUpdate_5[3:0]) begin
              TBEMemory_3_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_3_fields_0 <= _GEN_2492;
            end
          end else begin
            TBEMemory_3_fields_0 <= _GEN_2492;
          end
        end else begin
          TBEMemory_3_fields_0 <= _GEN_2492;
        end
      end else begin
        TBEMemory_3_fields_0 <= _GEN_3006;
      end
    end else if (_T_243) begin
      if (4'h3 == idxUpdate_7[3:0]) begin
        TBEMemory_3_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h3 == idxAlloc[3:0]) begin
          TBEMemory_3_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_3_fields_0 <= _GEN_3006;
        end
      end else if (_T_221) begin
        if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_fields_0 <= 32'h0;
        end else begin
          TBEMemory_3_fields_0 <= _GEN_3006;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h3 == idxUpdate_6[3:0]) begin
            TBEMemory_3_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_3_fields_0 <= _GEN_3006;
          end
        end else begin
          TBEMemory_3_fields_0 <= _GEN_3006;
        end
      end else begin
        TBEMemory_3_fields_0 <= _GEN_3006;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'h3 == idxUpdate_7[3:0]) begin
          TBEMemory_3_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEMemory_3_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_3_fields_0 <= _GEN_3006;
          end
        end else if (_T_221) begin
          if (4'h3 == idxUpdate_6[3:0]) begin
            TBEMemory_3_fields_0 <= 32'h0;
          end else begin
            TBEMemory_3_fields_0 <= _GEN_3006;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'h3 == idxUpdate_6[3:0]) begin
              TBEMemory_3_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_3_fields_0 <= _GEN_3006;
            end
          end else begin
            TBEMemory_3_fields_0 <= _GEN_3006;
          end
        end else begin
          TBEMemory_3_fields_0 <= _GEN_3006;
        end
      end else if (isAlloc_6) begin
        if (4'h3 == idxAlloc[3:0]) begin
          TBEMemory_3_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_3_fields_0 <= _GEN_3006;
        end
      end else if (_T_221) begin
        if (4'h3 == idxUpdate_6[3:0]) begin
          TBEMemory_3_fields_0 <= 32'h0;
        end else begin
          TBEMemory_3_fields_0 <= _GEN_3006;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h3 == idxUpdate_6[3:0]) begin
            TBEMemory_3_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_3_fields_0 <= _GEN_3006;
          end
        end else begin
          TBEMemory_3_fields_0 <= _GEN_3006;
        end
      end else begin
        TBEMemory_3_fields_0 <= _GEN_3006;
      end
    end else begin
      TBEMemory_3_fields_0 <= _GEN_3520;
    end
    if (reset) begin
      TBEMemory_4_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'h4 == idxAlloc[3:0]) begin
        TBEMemory_4_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h4 == idxAlloc[3:0]) begin
          TBEMemory_4_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEMemory_4_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEMemory_4_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEMemory_4_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEMemory_4_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEMemory_4_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEMemory_4_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEMemory_4_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h4 == idxUpdate_0[3:0]) begin
                        TBEMemory_4_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEMemory_4_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEMemory_4_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h4 == idxUpdate_0[3:0]) begin
                        TBEMemory_4_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h4 == idxAlloc[3:0]) begin
                        TBEMemory_4_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'h4 == idxUpdate_0[3:0]) begin
                        TBEMemory_4_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h4 == idxUpdate_0[3:0]) begin
                          TBEMemory_4_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEMemory_4_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEMemory_4_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h4 == idxUpdate_0[3:0]) begin
                        TBEMemory_4_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_4_state_state <= _GEN_469;
                end
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEMemory_4_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_4_state_state <= _GEN_469;
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_state_state <= 2'h0;
                  end else begin
                    TBEMemory_4_state_state <= _GEN_469;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_4_state_state <= _GEN_469;
                  end else if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_4_state_state <= _GEN_469;
                  end
                end else begin
                  TBEMemory_4_state_state <= _GEN_469;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEMemory_4_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_4_state_state <= _GEN_469;
                    end
                  end else if (_T_111) begin
                    if (4'h4 == idxUpdate_1[3:0]) begin
                      TBEMemory_4_state_state <= 2'h0;
                    end else begin
                      TBEMemory_4_state_state <= _GEN_469;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_4_state_state <= _GEN_469;
                    end else if (4'h4 == idxUpdate_1[3:0]) begin
                      TBEMemory_4_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_4_state_state <= _GEN_469;
                    end
                  end else begin
                    TBEMemory_4_state_state <= _GEN_469;
                  end
                end else if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEMemory_4_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_4_state_state <= _GEN_469;
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_state_state <= 2'h0;
                  end else begin
                    TBEMemory_4_state_state <= _GEN_469;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_4_state_state <= _GEN_469;
                  end else if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_4_state_state <= _GEN_469;
                  end
                end else begin
                  TBEMemory_4_state_state <= _GEN_469;
                end
              end else begin
                TBEMemory_4_state_state <= _GEN_983;
              end
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEMemory_4_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_4_state_state <= _GEN_983;
                end
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_state_state <= 2'h0;
                end else begin
                  TBEMemory_4_state_state <= _GEN_983;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_4_state_state <= _GEN_983;
                end else if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_4_state_state <= _GEN_983;
                end
              end else begin
                TBEMemory_4_state_state <= _GEN_983;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEMemory_4_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_4_state_state <= _GEN_983;
                  end
                end else if (_T_133) begin
                  if (4'h4 == idxUpdate_2[3:0]) begin
                    TBEMemory_4_state_state <= 2'h0;
                  end else begin
                    TBEMemory_4_state_state <= _GEN_983;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_4_state_state <= _GEN_983;
                  end else if (4'h4 == idxUpdate_2[3:0]) begin
                    TBEMemory_4_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_4_state_state <= _GEN_983;
                  end
                end else begin
                  TBEMemory_4_state_state <= _GEN_983;
                end
              end else if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEMemory_4_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_4_state_state <= _GEN_983;
                end
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_state_state <= 2'h0;
                end else begin
                  TBEMemory_4_state_state <= _GEN_983;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_4_state_state <= _GEN_983;
                end else if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_4_state_state <= _GEN_983;
                end
              end else begin
                TBEMemory_4_state_state <= _GEN_983;
              end
            end else begin
              TBEMemory_4_state_state <= _GEN_1497;
            end
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEMemory_4_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_4_state_state <= _GEN_1497;
              end
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_state_state <= 2'h0;
              end else begin
                TBEMemory_4_state_state <= _GEN_1497;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_4_state_state <= _GEN_1497;
              end else if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_4_state_state <= _GEN_1497;
              end
            end else begin
              TBEMemory_4_state_state <= _GEN_1497;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEMemory_4_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_4_state_state <= _GEN_1497;
                end
              end else if (_T_155) begin
                if (4'h4 == idxUpdate_3[3:0]) begin
                  TBEMemory_4_state_state <= 2'h0;
                end else begin
                  TBEMemory_4_state_state <= _GEN_1497;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_4_state_state <= _GEN_1497;
                end else if (4'h4 == idxUpdate_3[3:0]) begin
                  TBEMemory_4_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_4_state_state <= _GEN_1497;
                end
              end else begin
                TBEMemory_4_state_state <= _GEN_1497;
              end
            end else if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEMemory_4_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_4_state_state <= _GEN_1497;
              end
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_state_state <= 2'h0;
              end else begin
                TBEMemory_4_state_state <= _GEN_1497;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_4_state_state <= _GEN_1497;
              end else if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_4_state_state <= _GEN_1497;
              end
            end else begin
              TBEMemory_4_state_state <= _GEN_1497;
            end
          end else begin
            TBEMemory_4_state_state <= _GEN_2011;
          end
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEMemory_4_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_4_state_state <= _GEN_2011;
            end
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_state_state <= 2'h0;
            end else begin
              TBEMemory_4_state_state <= _GEN_2011;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_4_state_state <= _GEN_2011;
            end else if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_4_state_state <= _GEN_2011;
            end
          end else begin
            TBEMemory_4_state_state <= _GEN_2011;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEMemory_4_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_4_state_state <= _GEN_2011;
              end
            end else if (_T_177) begin
              if (4'h4 == idxUpdate_4[3:0]) begin
                TBEMemory_4_state_state <= 2'h0;
              end else begin
                TBEMemory_4_state_state <= _GEN_2011;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_4_state_state <= _GEN_2011;
              end else if (4'h4 == idxUpdate_4[3:0]) begin
                TBEMemory_4_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_4_state_state <= _GEN_2011;
              end
            end else begin
              TBEMemory_4_state_state <= _GEN_2011;
            end
          end else if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEMemory_4_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_4_state_state <= _GEN_2011;
            end
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_state_state <= 2'h0;
            end else begin
              TBEMemory_4_state_state <= _GEN_2011;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_4_state_state <= _GEN_2011;
            end else if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_4_state_state <= _GEN_2011;
            end
          end else begin
            TBEMemory_4_state_state <= _GEN_2011;
          end
        end else begin
          TBEMemory_4_state_state <= _GEN_2525;
        end
      end else if (_T_221) begin
        if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEMemory_4_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_4_state_state <= _GEN_2525;
          end
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_state_state <= 2'h0;
          end else begin
            TBEMemory_4_state_state <= _GEN_2525;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_4_state_state <= _GEN_2525;
          end else if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_4_state_state <= _GEN_2525;
          end
        end else begin
          TBEMemory_4_state_state <= _GEN_2525;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEMemory_4_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_4_state_state <= _GEN_2525;
            end
          end else if (_T_199) begin
            if (4'h4 == idxUpdate_5[3:0]) begin
              TBEMemory_4_state_state <= 2'h0;
            end else begin
              TBEMemory_4_state_state <= _GEN_2525;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_4_state_state <= _GEN_2525;
            end else if (4'h4 == idxUpdate_5[3:0]) begin
              TBEMemory_4_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_4_state_state <= _GEN_2525;
            end
          end else begin
            TBEMemory_4_state_state <= _GEN_2525;
          end
        end else if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEMemory_4_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_4_state_state <= _GEN_2525;
          end
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_state_state <= 2'h0;
          end else begin
            TBEMemory_4_state_state <= _GEN_2525;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_4_state_state <= _GEN_2525;
          end else if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_4_state_state <= _GEN_2525;
          end
        end else begin
          TBEMemory_4_state_state <= _GEN_2525;
        end
      end else begin
        TBEMemory_4_state_state <= _GEN_3039;
      end
    end else if (_T_243) begin
      if (4'h4 == idxUpdate_7[3:0]) begin
        TBEMemory_4_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'h4 == idxAlloc[3:0]) begin
          TBEMemory_4_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_4_state_state <= _GEN_3039;
        end
      end else if (_T_221) begin
        if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_state_state <= 2'h0;
        end else begin
          TBEMemory_4_state_state <= _GEN_3039;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_4_state_state <= _GEN_3039;
        end else if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_4_state_state <= _GEN_3039;
        end
      end else begin
        TBEMemory_4_state_state <= _GEN_3039;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEMemory_4_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_4_state_state <= _GEN_3039;
          end
        end else if (_T_221) begin
          if (4'h4 == idxUpdate_6[3:0]) begin
            TBEMemory_4_state_state <= 2'h0;
          end else begin
            TBEMemory_4_state_state <= _GEN_3039;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_4_state_state <= _GEN_3039;
          end else if (4'h4 == idxUpdate_6[3:0]) begin
            TBEMemory_4_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_4_state_state <= _GEN_3039;
          end
        end else begin
          TBEMemory_4_state_state <= _GEN_3039;
        end
      end else if (4'h4 == idxUpdate_7[3:0]) begin
        TBEMemory_4_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h4 == idxAlloc[3:0]) begin
          TBEMemory_4_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_4_state_state <= _GEN_3039;
        end
      end else if (_T_221) begin
        if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_state_state <= 2'h0;
        end else begin
          TBEMemory_4_state_state <= _GEN_3039;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_4_state_state <= _GEN_3039;
        end else if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_4_state_state <= _GEN_3039;
        end
      end else begin
        TBEMemory_4_state_state <= _GEN_3039;
      end
    end else begin
      TBEMemory_4_state_state <= _GEN_3553;
    end
    if (reset) begin
      TBEMemory_4_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'h4 == idxAlloc[3:0]) begin
        TBEMemory_4_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h4 == idxAlloc[3:0]) begin
          TBEMemory_4_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEMemory_4_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEMemory_4_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEMemory_4_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEMemory_4_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEMemory_4_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEMemory_4_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEMemory_4_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h4 == idxUpdate_0[3:0]) begin
                        TBEMemory_4_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEMemory_4_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEMemory_4_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h4 == idxUpdate_0[3:0]) begin
                        TBEMemory_4_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h4 == idxAlloc[3:0]) begin
                        TBEMemory_4_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'h4 == idxUpdate_0[3:0]) begin
                        TBEMemory_4_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h4 == idxUpdate_0[3:0]) begin
                          TBEMemory_4_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEMemory_4_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEMemory_4_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h4 == idxUpdate_0[3:0]) begin
                        TBEMemory_4_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_4_way <= _GEN_453;
                end
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEMemory_4_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_4_way <= _GEN_453;
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_way <= 3'h2;
                  end else begin
                    TBEMemory_4_way <= _GEN_453;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_4_way <= _GEN_453;
                  end else if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_4_way <= _GEN_453;
                  end
                end else begin
                  TBEMemory_4_way <= _GEN_453;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEMemory_4_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_4_way <= _GEN_453;
                    end
                  end else if (_T_111) begin
                    if (4'h4 == idxUpdate_1[3:0]) begin
                      TBEMemory_4_way <= 3'h2;
                    end else begin
                      TBEMemory_4_way <= _GEN_453;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_4_way <= _GEN_453;
                    end else if (4'h4 == idxUpdate_1[3:0]) begin
                      TBEMemory_4_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_4_way <= _GEN_453;
                    end
                  end else begin
                    TBEMemory_4_way <= _GEN_453;
                  end
                end else if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEMemory_4_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_4_way <= _GEN_453;
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_way <= 3'h2;
                  end else begin
                    TBEMemory_4_way <= _GEN_453;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_4_way <= _GEN_453;
                  end else if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_4_way <= _GEN_453;
                  end
                end else begin
                  TBEMemory_4_way <= _GEN_453;
                end
              end else begin
                TBEMemory_4_way <= _GEN_967;
              end
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEMemory_4_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_4_way <= _GEN_967;
                end
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_way <= 3'h2;
                end else begin
                  TBEMemory_4_way <= _GEN_967;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_4_way <= _GEN_967;
                end else if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_4_way <= _GEN_967;
                end
              end else begin
                TBEMemory_4_way <= _GEN_967;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEMemory_4_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_4_way <= _GEN_967;
                  end
                end else if (_T_133) begin
                  if (4'h4 == idxUpdate_2[3:0]) begin
                    TBEMemory_4_way <= 3'h2;
                  end else begin
                    TBEMemory_4_way <= _GEN_967;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_4_way <= _GEN_967;
                  end else if (4'h4 == idxUpdate_2[3:0]) begin
                    TBEMemory_4_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_4_way <= _GEN_967;
                  end
                end else begin
                  TBEMemory_4_way <= _GEN_967;
                end
              end else if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEMemory_4_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_4_way <= _GEN_967;
                end
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_way <= 3'h2;
                end else begin
                  TBEMemory_4_way <= _GEN_967;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_4_way <= _GEN_967;
                end else if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_4_way <= _GEN_967;
                end
              end else begin
                TBEMemory_4_way <= _GEN_967;
              end
            end else begin
              TBEMemory_4_way <= _GEN_1481;
            end
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEMemory_4_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_4_way <= _GEN_1481;
              end
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_way <= 3'h2;
              end else begin
                TBEMemory_4_way <= _GEN_1481;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_4_way <= _GEN_1481;
              end else if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_4_way <= _GEN_1481;
              end
            end else begin
              TBEMemory_4_way <= _GEN_1481;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEMemory_4_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_4_way <= _GEN_1481;
                end
              end else if (_T_155) begin
                if (4'h4 == idxUpdate_3[3:0]) begin
                  TBEMemory_4_way <= 3'h2;
                end else begin
                  TBEMemory_4_way <= _GEN_1481;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_4_way <= _GEN_1481;
                end else if (4'h4 == idxUpdate_3[3:0]) begin
                  TBEMemory_4_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_4_way <= _GEN_1481;
                end
              end else begin
                TBEMemory_4_way <= _GEN_1481;
              end
            end else if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEMemory_4_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_4_way <= _GEN_1481;
              end
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_way <= 3'h2;
              end else begin
                TBEMemory_4_way <= _GEN_1481;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_4_way <= _GEN_1481;
              end else if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_4_way <= _GEN_1481;
              end
            end else begin
              TBEMemory_4_way <= _GEN_1481;
            end
          end else begin
            TBEMemory_4_way <= _GEN_1995;
          end
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEMemory_4_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_4_way <= _GEN_1995;
            end
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_way <= 3'h2;
            end else begin
              TBEMemory_4_way <= _GEN_1995;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_4_way <= _GEN_1995;
            end else if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_4_way <= _GEN_1995;
            end
          end else begin
            TBEMemory_4_way <= _GEN_1995;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEMemory_4_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_4_way <= _GEN_1995;
              end
            end else if (_T_177) begin
              if (4'h4 == idxUpdate_4[3:0]) begin
                TBEMemory_4_way <= 3'h2;
              end else begin
                TBEMemory_4_way <= _GEN_1995;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_4_way <= _GEN_1995;
              end else if (4'h4 == idxUpdate_4[3:0]) begin
                TBEMemory_4_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_4_way <= _GEN_1995;
              end
            end else begin
              TBEMemory_4_way <= _GEN_1995;
            end
          end else if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEMemory_4_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_4_way <= _GEN_1995;
            end
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_way <= 3'h2;
            end else begin
              TBEMemory_4_way <= _GEN_1995;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_4_way <= _GEN_1995;
            end else if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_4_way <= _GEN_1995;
            end
          end else begin
            TBEMemory_4_way <= _GEN_1995;
          end
        end else begin
          TBEMemory_4_way <= _GEN_2509;
        end
      end else if (_T_221) begin
        if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEMemory_4_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_4_way <= _GEN_2509;
          end
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_way <= 3'h2;
          end else begin
            TBEMemory_4_way <= _GEN_2509;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_4_way <= _GEN_2509;
          end else if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_4_way <= _GEN_2509;
          end
        end else begin
          TBEMemory_4_way <= _GEN_2509;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEMemory_4_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_4_way <= _GEN_2509;
            end
          end else if (_T_199) begin
            if (4'h4 == idxUpdate_5[3:0]) begin
              TBEMemory_4_way <= 3'h2;
            end else begin
              TBEMemory_4_way <= _GEN_2509;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_4_way <= _GEN_2509;
            end else if (4'h4 == idxUpdate_5[3:0]) begin
              TBEMemory_4_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_4_way <= _GEN_2509;
            end
          end else begin
            TBEMemory_4_way <= _GEN_2509;
          end
        end else if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEMemory_4_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_4_way <= _GEN_2509;
          end
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_way <= 3'h2;
          end else begin
            TBEMemory_4_way <= _GEN_2509;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_4_way <= _GEN_2509;
          end else if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_4_way <= _GEN_2509;
          end
        end else begin
          TBEMemory_4_way <= _GEN_2509;
        end
      end else begin
        TBEMemory_4_way <= _GEN_3023;
      end
    end else if (_T_243) begin
      if (4'h4 == idxUpdate_7[3:0]) begin
        TBEMemory_4_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'h4 == idxAlloc[3:0]) begin
          TBEMemory_4_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_4_way <= _GEN_3023;
        end
      end else if (_T_221) begin
        if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_way <= 3'h2;
        end else begin
          TBEMemory_4_way <= _GEN_3023;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_4_way <= _GEN_3023;
        end else if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_4_way <= _GEN_3023;
        end
      end else begin
        TBEMemory_4_way <= _GEN_3023;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEMemory_4_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_4_way <= _GEN_3023;
          end
        end else if (_T_221) begin
          if (4'h4 == idxUpdate_6[3:0]) begin
            TBEMemory_4_way <= 3'h2;
          end else begin
            TBEMemory_4_way <= _GEN_3023;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_4_way <= _GEN_3023;
          end else if (4'h4 == idxUpdate_6[3:0]) begin
            TBEMemory_4_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_4_way <= _GEN_3023;
          end
        end else begin
          TBEMemory_4_way <= _GEN_3023;
        end
      end else if (4'h4 == idxUpdate_7[3:0]) begin
        TBEMemory_4_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h4 == idxAlloc[3:0]) begin
          TBEMemory_4_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_4_way <= _GEN_3023;
        end
      end else if (_T_221) begin
        if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_way <= 3'h2;
        end else begin
          TBEMemory_4_way <= _GEN_3023;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_4_way <= _GEN_3023;
        end else if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_4_way <= _GEN_3023;
        end
      end else begin
        TBEMemory_4_way <= _GEN_3023;
      end
    end else begin
      TBEMemory_4_way <= _GEN_3537;
    end
    if (reset) begin
      TBEMemory_4_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h4 == idxAlloc[3:0]) begin
        TBEMemory_4_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'h4 == idxAlloc[3:0]) begin
          TBEMemory_4_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEMemory_4_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEMemory_4_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEMemory_4_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEMemory_4_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEMemory_4_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEMemory_4_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEMemory_4_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h4 == idxUpdate_0[3:0]) begin
                        TBEMemory_4_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEMemory_4_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEMemory_4_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h4 == idxUpdate_0[3:0]) begin
                        TBEMemory_4_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h4 == idxUpdate_1[3:0]) begin
                      TBEMemory_4_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'h4 == idxAlloc[3:0]) begin
                        TBEMemory_4_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'h4 == idxUpdate_0[3:0]) begin
                        TBEMemory_4_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'h4 == idxUpdate_0[3:0]) begin
                          TBEMemory_4_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEMemory_4_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEMemory_4_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h4 == idxUpdate_0[3:0]) begin
                        TBEMemory_4_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_437;
                end
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEMemory_4_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_437;
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_437;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h4 == idxUpdate_1[3:0]) begin
                      TBEMemory_4_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_4_fields_0 <= _GEN_437;
                    end
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_437;
                  end
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_437;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h4 == idxUpdate_2[3:0]) begin
                    TBEMemory_4_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEMemory_4_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_4_fields_0 <= _GEN_437;
                    end
                  end else if (_T_111) begin
                    if (4'h4 == idxUpdate_1[3:0]) begin
                      TBEMemory_4_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_4_fields_0 <= _GEN_437;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'h4 == idxUpdate_1[3:0]) begin
                        TBEMemory_4_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_4_fields_0 <= _GEN_437;
                      end
                    end else begin
                      TBEMemory_4_fields_0 <= _GEN_437;
                    end
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_437;
                  end
                end else if (isAlloc_1) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEMemory_4_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_437;
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEMemory_4_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_437;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h4 == idxUpdate_1[3:0]) begin
                      TBEMemory_4_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_4_fields_0 <= _GEN_437;
                    end
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_437;
                  end
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_437;
                end
              end else begin
                TBEMemory_4_fields_0 <= _GEN_951;
              end
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEMemory_4_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_951;
                end
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_951;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h4 == idxUpdate_2[3:0]) begin
                    TBEMemory_4_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_951;
                  end
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_951;
                end
              end else begin
                TBEMemory_4_fields_0 <= _GEN_951;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h4 == idxUpdate_3[3:0]) begin
                  TBEMemory_4_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEMemory_4_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_951;
                  end
                end else if (_T_133) begin
                  if (4'h4 == idxUpdate_2[3:0]) begin
                    TBEMemory_4_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_951;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'h4 == idxUpdate_2[3:0]) begin
                      TBEMemory_4_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_4_fields_0 <= _GEN_951;
                    end
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_951;
                  end
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_951;
                end
              end else if (isAlloc_2) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEMemory_4_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_951;
                end
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEMemory_4_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_951;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h4 == idxUpdate_2[3:0]) begin
                    TBEMemory_4_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_951;
                  end
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_951;
                end
              end else begin
                TBEMemory_4_fields_0 <= _GEN_951;
              end
            end else begin
              TBEMemory_4_fields_0 <= _GEN_1465;
            end
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEMemory_4_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_4_fields_0 <= _GEN_1465;
              end
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_fields_0 <= 32'h0;
              end else begin
                TBEMemory_4_fields_0 <= _GEN_1465;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h4 == idxUpdate_3[3:0]) begin
                  TBEMemory_4_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_1465;
                end
              end else begin
                TBEMemory_4_fields_0 <= _GEN_1465;
              end
            end else begin
              TBEMemory_4_fields_0 <= _GEN_1465;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h4 == idxUpdate_4[3:0]) begin
                TBEMemory_4_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEMemory_4_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_1465;
                end
              end else if (_T_155) begin
                if (4'h4 == idxUpdate_3[3:0]) begin
                  TBEMemory_4_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_1465;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'h4 == idxUpdate_3[3:0]) begin
                    TBEMemory_4_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_4_fields_0 <= _GEN_1465;
                  end
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_1465;
                end
              end else begin
                TBEMemory_4_fields_0 <= _GEN_1465;
              end
            end else if (isAlloc_3) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEMemory_4_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_4_fields_0 <= _GEN_1465;
              end
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEMemory_4_fields_0 <= 32'h0;
              end else begin
                TBEMemory_4_fields_0 <= _GEN_1465;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h4 == idxUpdate_3[3:0]) begin
                  TBEMemory_4_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_1465;
                end
              end else begin
                TBEMemory_4_fields_0 <= _GEN_1465;
              end
            end else begin
              TBEMemory_4_fields_0 <= _GEN_1465;
            end
          end else begin
            TBEMemory_4_fields_0 <= _GEN_1979;
          end
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEMemory_4_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_4_fields_0 <= _GEN_1979;
            end
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_fields_0 <= 32'h0;
            end else begin
              TBEMemory_4_fields_0 <= _GEN_1979;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h4 == idxUpdate_4[3:0]) begin
                TBEMemory_4_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_4_fields_0 <= _GEN_1979;
              end
            end else begin
              TBEMemory_4_fields_0 <= _GEN_1979;
            end
          end else begin
            TBEMemory_4_fields_0 <= _GEN_1979;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h4 == idxUpdate_5[3:0]) begin
              TBEMemory_4_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEMemory_4_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_4_fields_0 <= _GEN_1979;
              end
            end else if (_T_177) begin
              if (4'h4 == idxUpdate_4[3:0]) begin
                TBEMemory_4_fields_0 <= 32'h0;
              end else begin
                TBEMemory_4_fields_0 <= _GEN_1979;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'h4 == idxUpdate_4[3:0]) begin
                  TBEMemory_4_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_4_fields_0 <= _GEN_1979;
                end
              end else begin
                TBEMemory_4_fields_0 <= _GEN_1979;
              end
            end else begin
              TBEMemory_4_fields_0 <= _GEN_1979;
            end
          end else if (isAlloc_4) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEMemory_4_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_4_fields_0 <= _GEN_1979;
            end
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEMemory_4_fields_0 <= 32'h0;
            end else begin
              TBEMemory_4_fields_0 <= _GEN_1979;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h4 == idxUpdate_4[3:0]) begin
                TBEMemory_4_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_4_fields_0 <= _GEN_1979;
              end
            end else begin
              TBEMemory_4_fields_0 <= _GEN_1979;
            end
          end else begin
            TBEMemory_4_fields_0 <= _GEN_1979;
          end
        end else begin
          TBEMemory_4_fields_0 <= _GEN_2493;
        end
      end else if (_T_221) begin
        if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEMemory_4_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_4_fields_0 <= _GEN_2493;
          end
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_fields_0 <= 32'h0;
          end else begin
            TBEMemory_4_fields_0 <= _GEN_2493;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h4 == idxUpdate_5[3:0]) begin
              TBEMemory_4_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_4_fields_0 <= _GEN_2493;
            end
          end else begin
            TBEMemory_4_fields_0 <= _GEN_2493;
          end
        end else begin
          TBEMemory_4_fields_0 <= _GEN_2493;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h4 == idxUpdate_6[3:0]) begin
            TBEMemory_4_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEMemory_4_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_4_fields_0 <= _GEN_2493;
            end
          end else if (_T_199) begin
            if (4'h4 == idxUpdate_5[3:0]) begin
              TBEMemory_4_fields_0 <= 32'h0;
            end else begin
              TBEMemory_4_fields_0 <= _GEN_2493;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'h4 == idxUpdate_5[3:0]) begin
                TBEMemory_4_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_4_fields_0 <= _GEN_2493;
              end
            end else begin
              TBEMemory_4_fields_0 <= _GEN_2493;
            end
          end else begin
            TBEMemory_4_fields_0 <= _GEN_2493;
          end
        end else if (isAlloc_5) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEMemory_4_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_4_fields_0 <= _GEN_2493;
          end
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEMemory_4_fields_0 <= 32'h0;
          end else begin
            TBEMemory_4_fields_0 <= _GEN_2493;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h4 == idxUpdate_5[3:0]) begin
              TBEMemory_4_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_4_fields_0 <= _GEN_2493;
            end
          end else begin
            TBEMemory_4_fields_0 <= _GEN_2493;
          end
        end else begin
          TBEMemory_4_fields_0 <= _GEN_2493;
        end
      end else begin
        TBEMemory_4_fields_0 <= _GEN_3007;
      end
    end else if (_T_243) begin
      if (4'h4 == idxUpdate_7[3:0]) begin
        TBEMemory_4_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h4 == idxAlloc[3:0]) begin
          TBEMemory_4_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_4_fields_0 <= _GEN_3007;
        end
      end else if (_T_221) begin
        if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_fields_0 <= 32'h0;
        end else begin
          TBEMemory_4_fields_0 <= _GEN_3007;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h4 == idxUpdate_6[3:0]) begin
            TBEMemory_4_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_4_fields_0 <= _GEN_3007;
          end
        end else begin
          TBEMemory_4_fields_0 <= _GEN_3007;
        end
      end else begin
        TBEMemory_4_fields_0 <= _GEN_3007;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'h4 == idxUpdate_7[3:0]) begin
          TBEMemory_4_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEMemory_4_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_4_fields_0 <= _GEN_3007;
          end
        end else if (_T_221) begin
          if (4'h4 == idxUpdate_6[3:0]) begin
            TBEMemory_4_fields_0 <= 32'h0;
          end else begin
            TBEMemory_4_fields_0 <= _GEN_3007;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'h4 == idxUpdate_6[3:0]) begin
              TBEMemory_4_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_4_fields_0 <= _GEN_3007;
            end
          end else begin
            TBEMemory_4_fields_0 <= _GEN_3007;
          end
        end else begin
          TBEMemory_4_fields_0 <= _GEN_3007;
        end
      end else if (isAlloc_6) begin
        if (4'h4 == idxAlloc[3:0]) begin
          TBEMemory_4_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_4_fields_0 <= _GEN_3007;
        end
      end else if (_T_221) begin
        if (4'h4 == idxUpdate_6[3:0]) begin
          TBEMemory_4_fields_0 <= 32'h0;
        end else begin
          TBEMemory_4_fields_0 <= _GEN_3007;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h4 == idxUpdate_6[3:0]) begin
            TBEMemory_4_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_4_fields_0 <= _GEN_3007;
          end
        end else begin
          TBEMemory_4_fields_0 <= _GEN_3007;
        end
      end else begin
        TBEMemory_4_fields_0 <= _GEN_3007;
      end
    end else begin
      TBEMemory_4_fields_0 <= _GEN_3521;
    end
    if (reset) begin
      TBEMemory_5_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'h5 == idxAlloc[3:0]) begin
        TBEMemory_5_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h5 == idxAlloc[3:0]) begin
          TBEMemory_5_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEMemory_5_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEMemory_5_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEMemory_5_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEMemory_5_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEMemory_5_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEMemory_5_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEMemory_5_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h5 == idxUpdate_0[3:0]) begin
                        TBEMemory_5_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEMemory_5_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEMemory_5_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h5 == idxUpdate_0[3:0]) begin
                        TBEMemory_5_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h5 == idxAlloc[3:0]) begin
                        TBEMemory_5_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'h5 == idxUpdate_0[3:0]) begin
                        TBEMemory_5_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h5 == idxUpdate_0[3:0]) begin
                          TBEMemory_5_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEMemory_5_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEMemory_5_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h5 == idxUpdate_0[3:0]) begin
                        TBEMemory_5_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_5_state_state <= _GEN_470;
                end
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEMemory_5_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_5_state_state <= _GEN_470;
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_state_state <= 2'h0;
                  end else begin
                    TBEMemory_5_state_state <= _GEN_470;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_5_state_state <= _GEN_470;
                  end else if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_5_state_state <= _GEN_470;
                  end
                end else begin
                  TBEMemory_5_state_state <= _GEN_470;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEMemory_5_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_5_state_state <= _GEN_470;
                    end
                  end else if (_T_111) begin
                    if (4'h5 == idxUpdate_1[3:0]) begin
                      TBEMemory_5_state_state <= 2'h0;
                    end else begin
                      TBEMemory_5_state_state <= _GEN_470;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_5_state_state <= _GEN_470;
                    end else if (4'h5 == idxUpdate_1[3:0]) begin
                      TBEMemory_5_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_5_state_state <= _GEN_470;
                    end
                  end else begin
                    TBEMemory_5_state_state <= _GEN_470;
                  end
                end else if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEMemory_5_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_5_state_state <= _GEN_470;
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_state_state <= 2'h0;
                  end else begin
                    TBEMemory_5_state_state <= _GEN_470;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_5_state_state <= _GEN_470;
                  end else if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_5_state_state <= _GEN_470;
                  end
                end else begin
                  TBEMemory_5_state_state <= _GEN_470;
                end
              end else begin
                TBEMemory_5_state_state <= _GEN_984;
              end
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEMemory_5_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_5_state_state <= _GEN_984;
                end
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_state_state <= 2'h0;
                end else begin
                  TBEMemory_5_state_state <= _GEN_984;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_5_state_state <= _GEN_984;
                end else if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_5_state_state <= _GEN_984;
                end
              end else begin
                TBEMemory_5_state_state <= _GEN_984;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEMemory_5_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_5_state_state <= _GEN_984;
                  end
                end else if (_T_133) begin
                  if (4'h5 == idxUpdate_2[3:0]) begin
                    TBEMemory_5_state_state <= 2'h0;
                  end else begin
                    TBEMemory_5_state_state <= _GEN_984;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_5_state_state <= _GEN_984;
                  end else if (4'h5 == idxUpdate_2[3:0]) begin
                    TBEMemory_5_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_5_state_state <= _GEN_984;
                  end
                end else begin
                  TBEMemory_5_state_state <= _GEN_984;
                end
              end else if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEMemory_5_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_5_state_state <= _GEN_984;
                end
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_state_state <= 2'h0;
                end else begin
                  TBEMemory_5_state_state <= _GEN_984;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_5_state_state <= _GEN_984;
                end else if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_5_state_state <= _GEN_984;
                end
              end else begin
                TBEMemory_5_state_state <= _GEN_984;
              end
            end else begin
              TBEMemory_5_state_state <= _GEN_1498;
            end
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEMemory_5_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_5_state_state <= _GEN_1498;
              end
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_state_state <= 2'h0;
              end else begin
                TBEMemory_5_state_state <= _GEN_1498;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_5_state_state <= _GEN_1498;
              end else if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_5_state_state <= _GEN_1498;
              end
            end else begin
              TBEMemory_5_state_state <= _GEN_1498;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEMemory_5_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_5_state_state <= _GEN_1498;
                end
              end else if (_T_155) begin
                if (4'h5 == idxUpdate_3[3:0]) begin
                  TBEMemory_5_state_state <= 2'h0;
                end else begin
                  TBEMemory_5_state_state <= _GEN_1498;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_5_state_state <= _GEN_1498;
                end else if (4'h5 == idxUpdate_3[3:0]) begin
                  TBEMemory_5_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_5_state_state <= _GEN_1498;
                end
              end else begin
                TBEMemory_5_state_state <= _GEN_1498;
              end
            end else if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEMemory_5_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_5_state_state <= _GEN_1498;
              end
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_state_state <= 2'h0;
              end else begin
                TBEMemory_5_state_state <= _GEN_1498;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_5_state_state <= _GEN_1498;
              end else if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_5_state_state <= _GEN_1498;
              end
            end else begin
              TBEMemory_5_state_state <= _GEN_1498;
            end
          end else begin
            TBEMemory_5_state_state <= _GEN_2012;
          end
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEMemory_5_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_5_state_state <= _GEN_2012;
            end
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_state_state <= 2'h0;
            end else begin
              TBEMemory_5_state_state <= _GEN_2012;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_5_state_state <= _GEN_2012;
            end else if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_5_state_state <= _GEN_2012;
            end
          end else begin
            TBEMemory_5_state_state <= _GEN_2012;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEMemory_5_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_5_state_state <= _GEN_2012;
              end
            end else if (_T_177) begin
              if (4'h5 == idxUpdate_4[3:0]) begin
                TBEMemory_5_state_state <= 2'h0;
              end else begin
                TBEMemory_5_state_state <= _GEN_2012;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_5_state_state <= _GEN_2012;
              end else if (4'h5 == idxUpdate_4[3:0]) begin
                TBEMemory_5_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_5_state_state <= _GEN_2012;
              end
            end else begin
              TBEMemory_5_state_state <= _GEN_2012;
            end
          end else if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEMemory_5_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_5_state_state <= _GEN_2012;
            end
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_state_state <= 2'h0;
            end else begin
              TBEMemory_5_state_state <= _GEN_2012;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_5_state_state <= _GEN_2012;
            end else if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_5_state_state <= _GEN_2012;
            end
          end else begin
            TBEMemory_5_state_state <= _GEN_2012;
          end
        end else begin
          TBEMemory_5_state_state <= _GEN_2526;
        end
      end else if (_T_221) begin
        if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEMemory_5_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_5_state_state <= _GEN_2526;
          end
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_state_state <= 2'h0;
          end else begin
            TBEMemory_5_state_state <= _GEN_2526;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_5_state_state <= _GEN_2526;
          end else if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_5_state_state <= _GEN_2526;
          end
        end else begin
          TBEMemory_5_state_state <= _GEN_2526;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEMemory_5_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_5_state_state <= _GEN_2526;
            end
          end else if (_T_199) begin
            if (4'h5 == idxUpdate_5[3:0]) begin
              TBEMemory_5_state_state <= 2'h0;
            end else begin
              TBEMemory_5_state_state <= _GEN_2526;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_5_state_state <= _GEN_2526;
            end else if (4'h5 == idxUpdate_5[3:0]) begin
              TBEMemory_5_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_5_state_state <= _GEN_2526;
            end
          end else begin
            TBEMemory_5_state_state <= _GEN_2526;
          end
        end else if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEMemory_5_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_5_state_state <= _GEN_2526;
          end
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_state_state <= 2'h0;
          end else begin
            TBEMemory_5_state_state <= _GEN_2526;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_5_state_state <= _GEN_2526;
          end else if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_5_state_state <= _GEN_2526;
          end
        end else begin
          TBEMemory_5_state_state <= _GEN_2526;
        end
      end else begin
        TBEMemory_5_state_state <= _GEN_3040;
      end
    end else if (_T_243) begin
      if (4'h5 == idxUpdate_7[3:0]) begin
        TBEMemory_5_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'h5 == idxAlloc[3:0]) begin
          TBEMemory_5_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_5_state_state <= _GEN_3040;
        end
      end else if (_T_221) begin
        if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_state_state <= 2'h0;
        end else begin
          TBEMemory_5_state_state <= _GEN_3040;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_5_state_state <= _GEN_3040;
        end else if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_5_state_state <= _GEN_3040;
        end
      end else begin
        TBEMemory_5_state_state <= _GEN_3040;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEMemory_5_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_5_state_state <= _GEN_3040;
          end
        end else if (_T_221) begin
          if (4'h5 == idxUpdate_6[3:0]) begin
            TBEMemory_5_state_state <= 2'h0;
          end else begin
            TBEMemory_5_state_state <= _GEN_3040;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_5_state_state <= _GEN_3040;
          end else if (4'h5 == idxUpdate_6[3:0]) begin
            TBEMemory_5_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_5_state_state <= _GEN_3040;
          end
        end else begin
          TBEMemory_5_state_state <= _GEN_3040;
        end
      end else if (4'h5 == idxUpdate_7[3:0]) begin
        TBEMemory_5_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h5 == idxAlloc[3:0]) begin
          TBEMemory_5_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_5_state_state <= _GEN_3040;
        end
      end else if (_T_221) begin
        if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_state_state <= 2'h0;
        end else begin
          TBEMemory_5_state_state <= _GEN_3040;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_5_state_state <= _GEN_3040;
        end else if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_5_state_state <= _GEN_3040;
        end
      end else begin
        TBEMemory_5_state_state <= _GEN_3040;
      end
    end else begin
      TBEMemory_5_state_state <= _GEN_3554;
    end
    if (reset) begin
      TBEMemory_5_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'h5 == idxAlloc[3:0]) begin
        TBEMemory_5_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h5 == idxAlloc[3:0]) begin
          TBEMemory_5_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEMemory_5_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEMemory_5_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEMemory_5_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEMemory_5_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEMemory_5_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEMemory_5_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEMemory_5_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h5 == idxUpdate_0[3:0]) begin
                        TBEMemory_5_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEMemory_5_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEMemory_5_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h5 == idxUpdate_0[3:0]) begin
                        TBEMemory_5_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h5 == idxAlloc[3:0]) begin
                        TBEMemory_5_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'h5 == idxUpdate_0[3:0]) begin
                        TBEMemory_5_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h5 == idxUpdate_0[3:0]) begin
                          TBEMemory_5_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEMemory_5_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEMemory_5_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h5 == idxUpdate_0[3:0]) begin
                        TBEMemory_5_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_5_way <= _GEN_454;
                end
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEMemory_5_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_5_way <= _GEN_454;
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_way <= 3'h2;
                  end else begin
                    TBEMemory_5_way <= _GEN_454;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_5_way <= _GEN_454;
                  end else if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_5_way <= _GEN_454;
                  end
                end else begin
                  TBEMemory_5_way <= _GEN_454;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEMemory_5_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_5_way <= _GEN_454;
                    end
                  end else if (_T_111) begin
                    if (4'h5 == idxUpdate_1[3:0]) begin
                      TBEMemory_5_way <= 3'h2;
                    end else begin
                      TBEMemory_5_way <= _GEN_454;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_5_way <= _GEN_454;
                    end else if (4'h5 == idxUpdate_1[3:0]) begin
                      TBEMemory_5_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_5_way <= _GEN_454;
                    end
                  end else begin
                    TBEMemory_5_way <= _GEN_454;
                  end
                end else if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEMemory_5_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_5_way <= _GEN_454;
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_way <= 3'h2;
                  end else begin
                    TBEMemory_5_way <= _GEN_454;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_5_way <= _GEN_454;
                  end else if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_5_way <= _GEN_454;
                  end
                end else begin
                  TBEMemory_5_way <= _GEN_454;
                end
              end else begin
                TBEMemory_5_way <= _GEN_968;
              end
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEMemory_5_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_5_way <= _GEN_968;
                end
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_way <= 3'h2;
                end else begin
                  TBEMemory_5_way <= _GEN_968;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_5_way <= _GEN_968;
                end else if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_5_way <= _GEN_968;
                end
              end else begin
                TBEMemory_5_way <= _GEN_968;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEMemory_5_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_5_way <= _GEN_968;
                  end
                end else if (_T_133) begin
                  if (4'h5 == idxUpdate_2[3:0]) begin
                    TBEMemory_5_way <= 3'h2;
                  end else begin
                    TBEMemory_5_way <= _GEN_968;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_5_way <= _GEN_968;
                  end else if (4'h5 == idxUpdate_2[3:0]) begin
                    TBEMemory_5_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_5_way <= _GEN_968;
                  end
                end else begin
                  TBEMemory_5_way <= _GEN_968;
                end
              end else if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEMemory_5_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_5_way <= _GEN_968;
                end
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_way <= 3'h2;
                end else begin
                  TBEMemory_5_way <= _GEN_968;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_5_way <= _GEN_968;
                end else if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_5_way <= _GEN_968;
                end
              end else begin
                TBEMemory_5_way <= _GEN_968;
              end
            end else begin
              TBEMemory_5_way <= _GEN_1482;
            end
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEMemory_5_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_5_way <= _GEN_1482;
              end
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_way <= 3'h2;
              end else begin
                TBEMemory_5_way <= _GEN_1482;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_5_way <= _GEN_1482;
              end else if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_5_way <= _GEN_1482;
              end
            end else begin
              TBEMemory_5_way <= _GEN_1482;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEMemory_5_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_5_way <= _GEN_1482;
                end
              end else if (_T_155) begin
                if (4'h5 == idxUpdate_3[3:0]) begin
                  TBEMemory_5_way <= 3'h2;
                end else begin
                  TBEMemory_5_way <= _GEN_1482;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_5_way <= _GEN_1482;
                end else if (4'h5 == idxUpdate_3[3:0]) begin
                  TBEMemory_5_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_5_way <= _GEN_1482;
                end
              end else begin
                TBEMemory_5_way <= _GEN_1482;
              end
            end else if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEMemory_5_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_5_way <= _GEN_1482;
              end
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_way <= 3'h2;
              end else begin
                TBEMemory_5_way <= _GEN_1482;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_5_way <= _GEN_1482;
              end else if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_5_way <= _GEN_1482;
              end
            end else begin
              TBEMemory_5_way <= _GEN_1482;
            end
          end else begin
            TBEMemory_5_way <= _GEN_1996;
          end
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEMemory_5_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_5_way <= _GEN_1996;
            end
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_way <= 3'h2;
            end else begin
              TBEMemory_5_way <= _GEN_1996;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_5_way <= _GEN_1996;
            end else if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_5_way <= _GEN_1996;
            end
          end else begin
            TBEMemory_5_way <= _GEN_1996;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEMemory_5_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_5_way <= _GEN_1996;
              end
            end else if (_T_177) begin
              if (4'h5 == idxUpdate_4[3:0]) begin
                TBEMemory_5_way <= 3'h2;
              end else begin
                TBEMemory_5_way <= _GEN_1996;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_5_way <= _GEN_1996;
              end else if (4'h5 == idxUpdate_4[3:0]) begin
                TBEMemory_5_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_5_way <= _GEN_1996;
              end
            end else begin
              TBEMemory_5_way <= _GEN_1996;
            end
          end else if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEMemory_5_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_5_way <= _GEN_1996;
            end
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_way <= 3'h2;
            end else begin
              TBEMemory_5_way <= _GEN_1996;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_5_way <= _GEN_1996;
            end else if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_5_way <= _GEN_1996;
            end
          end else begin
            TBEMemory_5_way <= _GEN_1996;
          end
        end else begin
          TBEMemory_5_way <= _GEN_2510;
        end
      end else if (_T_221) begin
        if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEMemory_5_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_5_way <= _GEN_2510;
          end
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_way <= 3'h2;
          end else begin
            TBEMemory_5_way <= _GEN_2510;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_5_way <= _GEN_2510;
          end else if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_5_way <= _GEN_2510;
          end
        end else begin
          TBEMemory_5_way <= _GEN_2510;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEMemory_5_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_5_way <= _GEN_2510;
            end
          end else if (_T_199) begin
            if (4'h5 == idxUpdate_5[3:0]) begin
              TBEMemory_5_way <= 3'h2;
            end else begin
              TBEMemory_5_way <= _GEN_2510;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_5_way <= _GEN_2510;
            end else if (4'h5 == idxUpdate_5[3:0]) begin
              TBEMemory_5_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_5_way <= _GEN_2510;
            end
          end else begin
            TBEMemory_5_way <= _GEN_2510;
          end
        end else if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEMemory_5_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_5_way <= _GEN_2510;
          end
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_way <= 3'h2;
          end else begin
            TBEMemory_5_way <= _GEN_2510;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_5_way <= _GEN_2510;
          end else if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_5_way <= _GEN_2510;
          end
        end else begin
          TBEMemory_5_way <= _GEN_2510;
        end
      end else begin
        TBEMemory_5_way <= _GEN_3024;
      end
    end else if (_T_243) begin
      if (4'h5 == idxUpdate_7[3:0]) begin
        TBEMemory_5_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'h5 == idxAlloc[3:0]) begin
          TBEMemory_5_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_5_way <= _GEN_3024;
        end
      end else if (_T_221) begin
        if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_way <= 3'h2;
        end else begin
          TBEMemory_5_way <= _GEN_3024;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_5_way <= _GEN_3024;
        end else if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_5_way <= _GEN_3024;
        end
      end else begin
        TBEMemory_5_way <= _GEN_3024;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEMemory_5_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_5_way <= _GEN_3024;
          end
        end else if (_T_221) begin
          if (4'h5 == idxUpdate_6[3:0]) begin
            TBEMemory_5_way <= 3'h2;
          end else begin
            TBEMemory_5_way <= _GEN_3024;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_5_way <= _GEN_3024;
          end else if (4'h5 == idxUpdate_6[3:0]) begin
            TBEMemory_5_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_5_way <= _GEN_3024;
          end
        end else begin
          TBEMemory_5_way <= _GEN_3024;
        end
      end else if (4'h5 == idxUpdate_7[3:0]) begin
        TBEMemory_5_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h5 == idxAlloc[3:0]) begin
          TBEMemory_5_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_5_way <= _GEN_3024;
        end
      end else if (_T_221) begin
        if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_way <= 3'h2;
        end else begin
          TBEMemory_5_way <= _GEN_3024;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_5_way <= _GEN_3024;
        end else if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_5_way <= _GEN_3024;
        end
      end else begin
        TBEMemory_5_way <= _GEN_3024;
      end
    end else begin
      TBEMemory_5_way <= _GEN_3538;
    end
    if (reset) begin
      TBEMemory_5_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h5 == idxAlloc[3:0]) begin
        TBEMemory_5_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'h5 == idxAlloc[3:0]) begin
          TBEMemory_5_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEMemory_5_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEMemory_5_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEMemory_5_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEMemory_5_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEMemory_5_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEMemory_5_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEMemory_5_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h5 == idxUpdate_0[3:0]) begin
                        TBEMemory_5_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEMemory_5_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEMemory_5_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h5 == idxUpdate_0[3:0]) begin
                        TBEMemory_5_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h5 == idxUpdate_1[3:0]) begin
                      TBEMemory_5_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'h5 == idxAlloc[3:0]) begin
                        TBEMemory_5_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'h5 == idxUpdate_0[3:0]) begin
                        TBEMemory_5_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'h5 == idxUpdate_0[3:0]) begin
                          TBEMemory_5_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEMemory_5_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEMemory_5_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h5 == idxUpdate_0[3:0]) begin
                        TBEMemory_5_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_438;
                end
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEMemory_5_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_438;
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_438;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h5 == idxUpdate_1[3:0]) begin
                      TBEMemory_5_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_5_fields_0 <= _GEN_438;
                    end
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_438;
                  end
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_438;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h5 == idxUpdate_2[3:0]) begin
                    TBEMemory_5_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEMemory_5_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_5_fields_0 <= _GEN_438;
                    end
                  end else if (_T_111) begin
                    if (4'h5 == idxUpdate_1[3:0]) begin
                      TBEMemory_5_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_5_fields_0 <= _GEN_438;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'h5 == idxUpdate_1[3:0]) begin
                        TBEMemory_5_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_5_fields_0 <= _GEN_438;
                      end
                    end else begin
                      TBEMemory_5_fields_0 <= _GEN_438;
                    end
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_438;
                  end
                end else if (isAlloc_1) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEMemory_5_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_438;
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEMemory_5_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_438;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h5 == idxUpdate_1[3:0]) begin
                      TBEMemory_5_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_5_fields_0 <= _GEN_438;
                    end
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_438;
                  end
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_438;
                end
              end else begin
                TBEMemory_5_fields_0 <= _GEN_952;
              end
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEMemory_5_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_952;
                end
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_952;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h5 == idxUpdate_2[3:0]) begin
                    TBEMemory_5_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_952;
                  end
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_952;
                end
              end else begin
                TBEMemory_5_fields_0 <= _GEN_952;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h5 == idxUpdate_3[3:0]) begin
                  TBEMemory_5_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEMemory_5_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_952;
                  end
                end else if (_T_133) begin
                  if (4'h5 == idxUpdate_2[3:0]) begin
                    TBEMemory_5_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_952;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'h5 == idxUpdate_2[3:0]) begin
                      TBEMemory_5_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_5_fields_0 <= _GEN_952;
                    end
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_952;
                  end
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_952;
                end
              end else if (isAlloc_2) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEMemory_5_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_952;
                end
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEMemory_5_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_952;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h5 == idxUpdate_2[3:0]) begin
                    TBEMemory_5_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_952;
                  end
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_952;
                end
              end else begin
                TBEMemory_5_fields_0 <= _GEN_952;
              end
            end else begin
              TBEMemory_5_fields_0 <= _GEN_1466;
            end
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEMemory_5_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_5_fields_0 <= _GEN_1466;
              end
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_fields_0 <= 32'h0;
              end else begin
                TBEMemory_5_fields_0 <= _GEN_1466;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h5 == idxUpdate_3[3:0]) begin
                  TBEMemory_5_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_1466;
                end
              end else begin
                TBEMemory_5_fields_0 <= _GEN_1466;
              end
            end else begin
              TBEMemory_5_fields_0 <= _GEN_1466;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h5 == idxUpdate_4[3:0]) begin
                TBEMemory_5_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEMemory_5_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_1466;
                end
              end else if (_T_155) begin
                if (4'h5 == idxUpdate_3[3:0]) begin
                  TBEMemory_5_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_1466;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'h5 == idxUpdate_3[3:0]) begin
                    TBEMemory_5_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_5_fields_0 <= _GEN_1466;
                  end
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_1466;
                end
              end else begin
                TBEMemory_5_fields_0 <= _GEN_1466;
              end
            end else if (isAlloc_3) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEMemory_5_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_5_fields_0 <= _GEN_1466;
              end
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEMemory_5_fields_0 <= 32'h0;
              end else begin
                TBEMemory_5_fields_0 <= _GEN_1466;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h5 == idxUpdate_3[3:0]) begin
                  TBEMemory_5_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_1466;
                end
              end else begin
                TBEMemory_5_fields_0 <= _GEN_1466;
              end
            end else begin
              TBEMemory_5_fields_0 <= _GEN_1466;
            end
          end else begin
            TBEMemory_5_fields_0 <= _GEN_1980;
          end
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEMemory_5_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_5_fields_0 <= _GEN_1980;
            end
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_fields_0 <= 32'h0;
            end else begin
              TBEMemory_5_fields_0 <= _GEN_1980;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h5 == idxUpdate_4[3:0]) begin
                TBEMemory_5_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_5_fields_0 <= _GEN_1980;
              end
            end else begin
              TBEMemory_5_fields_0 <= _GEN_1980;
            end
          end else begin
            TBEMemory_5_fields_0 <= _GEN_1980;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h5 == idxUpdate_5[3:0]) begin
              TBEMemory_5_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEMemory_5_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_5_fields_0 <= _GEN_1980;
              end
            end else if (_T_177) begin
              if (4'h5 == idxUpdate_4[3:0]) begin
                TBEMemory_5_fields_0 <= 32'h0;
              end else begin
                TBEMemory_5_fields_0 <= _GEN_1980;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'h5 == idxUpdate_4[3:0]) begin
                  TBEMemory_5_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_5_fields_0 <= _GEN_1980;
                end
              end else begin
                TBEMemory_5_fields_0 <= _GEN_1980;
              end
            end else begin
              TBEMemory_5_fields_0 <= _GEN_1980;
            end
          end else if (isAlloc_4) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEMemory_5_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_5_fields_0 <= _GEN_1980;
            end
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEMemory_5_fields_0 <= 32'h0;
            end else begin
              TBEMemory_5_fields_0 <= _GEN_1980;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h5 == idxUpdate_4[3:0]) begin
                TBEMemory_5_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_5_fields_0 <= _GEN_1980;
              end
            end else begin
              TBEMemory_5_fields_0 <= _GEN_1980;
            end
          end else begin
            TBEMemory_5_fields_0 <= _GEN_1980;
          end
        end else begin
          TBEMemory_5_fields_0 <= _GEN_2494;
        end
      end else if (_T_221) begin
        if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEMemory_5_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_5_fields_0 <= _GEN_2494;
          end
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_fields_0 <= 32'h0;
          end else begin
            TBEMemory_5_fields_0 <= _GEN_2494;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h5 == idxUpdate_5[3:0]) begin
              TBEMemory_5_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_5_fields_0 <= _GEN_2494;
            end
          end else begin
            TBEMemory_5_fields_0 <= _GEN_2494;
          end
        end else begin
          TBEMemory_5_fields_0 <= _GEN_2494;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h5 == idxUpdate_6[3:0]) begin
            TBEMemory_5_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEMemory_5_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_5_fields_0 <= _GEN_2494;
            end
          end else if (_T_199) begin
            if (4'h5 == idxUpdate_5[3:0]) begin
              TBEMemory_5_fields_0 <= 32'h0;
            end else begin
              TBEMemory_5_fields_0 <= _GEN_2494;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'h5 == idxUpdate_5[3:0]) begin
                TBEMemory_5_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_5_fields_0 <= _GEN_2494;
              end
            end else begin
              TBEMemory_5_fields_0 <= _GEN_2494;
            end
          end else begin
            TBEMemory_5_fields_0 <= _GEN_2494;
          end
        end else if (isAlloc_5) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEMemory_5_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_5_fields_0 <= _GEN_2494;
          end
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEMemory_5_fields_0 <= 32'h0;
          end else begin
            TBEMemory_5_fields_0 <= _GEN_2494;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h5 == idxUpdate_5[3:0]) begin
              TBEMemory_5_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_5_fields_0 <= _GEN_2494;
            end
          end else begin
            TBEMemory_5_fields_0 <= _GEN_2494;
          end
        end else begin
          TBEMemory_5_fields_0 <= _GEN_2494;
        end
      end else begin
        TBEMemory_5_fields_0 <= _GEN_3008;
      end
    end else if (_T_243) begin
      if (4'h5 == idxUpdate_7[3:0]) begin
        TBEMemory_5_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h5 == idxAlloc[3:0]) begin
          TBEMemory_5_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_5_fields_0 <= _GEN_3008;
        end
      end else if (_T_221) begin
        if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_fields_0 <= 32'h0;
        end else begin
          TBEMemory_5_fields_0 <= _GEN_3008;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h5 == idxUpdate_6[3:0]) begin
            TBEMemory_5_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_5_fields_0 <= _GEN_3008;
          end
        end else begin
          TBEMemory_5_fields_0 <= _GEN_3008;
        end
      end else begin
        TBEMemory_5_fields_0 <= _GEN_3008;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'h5 == idxUpdate_7[3:0]) begin
          TBEMemory_5_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEMemory_5_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_5_fields_0 <= _GEN_3008;
          end
        end else if (_T_221) begin
          if (4'h5 == idxUpdate_6[3:0]) begin
            TBEMemory_5_fields_0 <= 32'h0;
          end else begin
            TBEMemory_5_fields_0 <= _GEN_3008;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'h5 == idxUpdate_6[3:0]) begin
              TBEMemory_5_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_5_fields_0 <= _GEN_3008;
            end
          end else begin
            TBEMemory_5_fields_0 <= _GEN_3008;
          end
        end else begin
          TBEMemory_5_fields_0 <= _GEN_3008;
        end
      end else if (isAlloc_6) begin
        if (4'h5 == idxAlloc[3:0]) begin
          TBEMemory_5_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_5_fields_0 <= _GEN_3008;
        end
      end else if (_T_221) begin
        if (4'h5 == idxUpdate_6[3:0]) begin
          TBEMemory_5_fields_0 <= 32'h0;
        end else begin
          TBEMemory_5_fields_0 <= _GEN_3008;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h5 == idxUpdate_6[3:0]) begin
            TBEMemory_5_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_5_fields_0 <= _GEN_3008;
          end
        end else begin
          TBEMemory_5_fields_0 <= _GEN_3008;
        end
      end else begin
        TBEMemory_5_fields_0 <= _GEN_3008;
      end
    end else begin
      TBEMemory_5_fields_0 <= _GEN_3522;
    end
    if (reset) begin
      TBEMemory_6_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'h6 == idxAlloc[3:0]) begin
        TBEMemory_6_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h6 == idxAlloc[3:0]) begin
          TBEMemory_6_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEMemory_6_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEMemory_6_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEMemory_6_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEMemory_6_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEMemory_6_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEMemory_6_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEMemory_6_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h6 == idxUpdate_0[3:0]) begin
                        TBEMemory_6_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEMemory_6_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEMemory_6_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h6 == idxUpdate_0[3:0]) begin
                        TBEMemory_6_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h6 == idxAlloc[3:0]) begin
                        TBEMemory_6_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'h6 == idxUpdate_0[3:0]) begin
                        TBEMemory_6_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h6 == idxUpdate_0[3:0]) begin
                          TBEMemory_6_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEMemory_6_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEMemory_6_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h6 == idxUpdate_0[3:0]) begin
                        TBEMemory_6_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_6_state_state <= _GEN_471;
                end
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEMemory_6_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_6_state_state <= _GEN_471;
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_state_state <= 2'h0;
                  end else begin
                    TBEMemory_6_state_state <= _GEN_471;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_6_state_state <= _GEN_471;
                  end else if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_6_state_state <= _GEN_471;
                  end
                end else begin
                  TBEMemory_6_state_state <= _GEN_471;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEMemory_6_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_6_state_state <= _GEN_471;
                    end
                  end else if (_T_111) begin
                    if (4'h6 == idxUpdate_1[3:0]) begin
                      TBEMemory_6_state_state <= 2'h0;
                    end else begin
                      TBEMemory_6_state_state <= _GEN_471;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_6_state_state <= _GEN_471;
                    end else if (4'h6 == idxUpdate_1[3:0]) begin
                      TBEMemory_6_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_6_state_state <= _GEN_471;
                    end
                  end else begin
                    TBEMemory_6_state_state <= _GEN_471;
                  end
                end else if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEMemory_6_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_6_state_state <= _GEN_471;
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_state_state <= 2'h0;
                  end else begin
                    TBEMemory_6_state_state <= _GEN_471;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_6_state_state <= _GEN_471;
                  end else if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_6_state_state <= _GEN_471;
                  end
                end else begin
                  TBEMemory_6_state_state <= _GEN_471;
                end
              end else begin
                TBEMemory_6_state_state <= _GEN_985;
              end
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEMemory_6_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_6_state_state <= _GEN_985;
                end
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_state_state <= 2'h0;
                end else begin
                  TBEMemory_6_state_state <= _GEN_985;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_6_state_state <= _GEN_985;
                end else if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_6_state_state <= _GEN_985;
                end
              end else begin
                TBEMemory_6_state_state <= _GEN_985;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEMemory_6_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_6_state_state <= _GEN_985;
                  end
                end else if (_T_133) begin
                  if (4'h6 == idxUpdate_2[3:0]) begin
                    TBEMemory_6_state_state <= 2'h0;
                  end else begin
                    TBEMemory_6_state_state <= _GEN_985;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_6_state_state <= _GEN_985;
                  end else if (4'h6 == idxUpdate_2[3:0]) begin
                    TBEMemory_6_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_6_state_state <= _GEN_985;
                  end
                end else begin
                  TBEMemory_6_state_state <= _GEN_985;
                end
              end else if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEMemory_6_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_6_state_state <= _GEN_985;
                end
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_state_state <= 2'h0;
                end else begin
                  TBEMemory_6_state_state <= _GEN_985;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_6_state_state <= _GEN_985;
                end else if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_6_state_state <= _GEN_985;
                end
              end else begin
                TBEMemory_6_state_state <= _GEN_985;
              end
            end else begin
              TBEMemory_6_state_state <= _GEN_1499;
            end
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEMemory_6_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_6_state_state <= _GEN_1499;
              end
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_state_state <= 2'h0;
              end else begin
                TBEMemory_6_state_state <= _GEN_1499;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_6_state_state <= _GEN_1499;
              end else if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_6_state_state <= _GEN_1499;
              end
            end else begin
              TBEMemory_6_state_state <= _GEN_1499;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEMemory_6_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_6_state_state <= _GEN_1499;
                end
              end else if (_T_155) begin
                if (4'h6 == idxUpdate_3[3:0]) begin
                  TBEMemory_6_state_state <= 2'h0;
                end else begin
                  TBEMemory_6_state_state <= _GEN_1499;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_6_state_state <= _GEN_1499;
                end else if (4'h6 == idxUpdate_3[3:0]) begin
                  TBEMemory_6_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_6_state_state <= _GEN_1499;
                end
              end else begin
                TBEMemory_6_state_state <= _GEN_1499;
              end
            end else if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEMemory_6_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_6_state_state <= _GEN_1499;
              end
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_state_state <= 2'h0;
              end else begin
                TBEMemory_6_state_state <= _GEN_1499;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_6_state_state <= _GEN_1499;
              end else if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_6_state_state <= _GEN_1499;
              end
            end else begin
              TBEMemory_6_state_state <= _GEN_1499;
            end
          end else begin
            TBEMemory_6_state_state <= _GEN_2013;
          end
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEMemory_6_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_6_state_state <= _GEN_2013;
            end
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_state_state <= 2'h0;
            end else begin
              TBEMemory_6_state_state <= _GEN_2013;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_6_state_state <= _GEN_2013;
            end else if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_6_state_state <= _GEN_2013;
            end
          end else begin
            TBEMemory_6_state_state <= _GEN_2013;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEMemory_6_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_6_state_state <= _GEN_2013;
              end
            end else if (_T_177) begin
              if (4'h6 == idxUpdate_4[3:0]) begin
                TBEMemory_6_state_state <= 2'h0;
              end else begin
                TBEMemory_6_state_state <= _GEN_2013;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_6_state_state <= _GEN_2013;
              end else if (4'h6 == idxUpdate_4[3:0]) begin
                TBEMemory_6_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_6_state_state <= _GEN_2013;
              end
            end else begin
              TBEMemory_6_state_state <= _GEN_2013;
            end
          end else if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEMemory_6_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_6_state_state <= _GEN_2013;
            end
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_state_state <= 2'h0;
            end else begin
              TBEMemory_6_state_state <= _GEN_2013;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_6_state_state <= _GEN_2013;
            end else if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_6_state_state <= _GEN_2013;
            end
          end else begin
            TBEMemory_6_state_state <= _GEN_2013;
          end
        end else begin
          TBEMemory_6_state_state <= _GEN_2527;
        end
      end else if (_T_221) begin
        if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEMemory_6_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_6_state_state <= _GEN_2527;
          end
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_state_state <= 2'h0;
          end else begin
            TBEMemory_6_state_state <= _GEN_2527;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_6_state_state <= _GEN_2527;
          end else if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_6_state_state <= _GEN_2527;
          end
        end else begin
          TBEMemory_6_state_state <= _GEN_2527;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEMemory_6_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_6_state_state <= _GEN_2527;
            end
          end else if (_T_199) begin
            if (4'h6 == idxUpdate_5[3:0]) begin
              TBEMemory_6_state_state <= 2'h0;
            end else begin
              TBEMemory_6_state_state <= _GEN_2527;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_6_state_state <= _GEN_2527;
            end else if (4'h6 == idxUpdate_5[3:0]) begin
              TBEMemory_6_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_6_state_state <= _GEN_2527;
            end
          end else begin
            TBEMemory_6_state_state <= _GEN_2527;
          end
        end else if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEMemory_6_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_6_state_state <= _GEN_2527;
          end
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_state_state <= 2'h0;
          end else begin
            TBEMemory_6_state_state <= _GEN_2527;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_6_state_state <= _GEN_2527;
          end else if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_6_state_state <= _GEN_2527;
          end
        end else begin
          TBEMemory_6_state_state <= _GEN_2527;
        end
      end else begin
        TBEMemory_6_state_state <= _GEN_3041;
      end
    end else if (_T_243) begin
      if (4'h6 == idxUpdate_7[3:0]) begin
        TBEMemory_6_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'h6 == idxAlloc[3:0]) begin
          TBEMemory_6_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_6_state_state <= _GEN_3041;
        end
      end else if (_T_221) begin
        if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_state_state <= 2'h0;
        end else begin
          TBEMemory_6_state_state <= _GEN_3041;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_6_state_state <= _GEN_3041;
        end else if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_6_state_state <= _GEN_3041;
        end
      end else begin
        TBEMemory_6_state_state <= _GEN_3041;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEMemory_6_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_6_state_state <= _GEN_3041;
          end
        end else if (_T_221) begin
          if (4'h6 == idxUpdate_6[3:0]) begin
            TBEMemory_6_state_state <= 2'h0;
          end else begin
            TBEMemory_6_state_state <= _GEN_3041;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_6_state_state <= _GEN_3041;
          end else if (4'h6 == idxUpdate_6[3:0]) begin
            TBEMemory_6_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_6_state_state <= _GEN_3041;
          end
        end else begin
          TBEMemory_6_state_state <= _GEN_3041;
        end
      end else if (4'h6 == idxUpdate_7[3:0]) begin
        TBEMemory_6_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h6 == idxAlloc[3:0]) begin
          TBEMemory_6_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_6_state_state <= _GEN_3041;
        end
      end else if (_T_221) begin
        if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_state_state <= 2'h0;
        end else begin
          TBEMemory_6_state_state <= _GEN_3041;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_6_state_state <= _GEN_3041;
        end else if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_6_state_state <= _GEN_3041;
        end
      end else begin
        TBEMemory_6_state_state <= _GEN_3041;
      end
    end else begin
      TBEMemory_6_state_state <= _GEN_3555;
    end
    if (reset) begin
      TBEMemory_6_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'h6 == idxAlloc[3:0]) begin
        TBEMemory_6_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h6 == idxAlloc[3:0]) begin
          TBEMemory_6_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEMemory_6_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEMemory_6_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEMemory_6_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEMemory_6_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEMemory_6_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEMemory_6_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEMemory_6_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h6 == idxUpdate_0[3:0]) begin
                        TBEMemory_6_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEMemory_6_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEMemory_6_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h6 == idxUpdate_0[3:0]) begin
                        TBEMemory_6_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h6 == idxAlloc[3:0]) begin
                        TBEMemory_6_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'h6 == idxUpdate_0[3:0]) begin
                        TBEMemory_6_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h6 == idxUpdate_0[3:0]) begin
                          TBEMemory_6_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEMemory_6_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEMemory_6_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h6 == idxUpdate_0[3:0]) begin
                        TBEMemory_6_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_6_way <= _GEN_455;
                end
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEMemory_6_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_6_way <= _GEN_455;
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_way <= 3'h2;
                  end else begin
                    TBEMemory_6_way <= _GEN_455;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_6_way <= _GEN_455;
                  end else if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_6_way <= _GEN_455;
                  end
                end else begin
                  TBEMemory_6_way <= _GEN_455;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEMemory_6_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_6_way <= _GEN_455;
                    end
                  end else if (_T_111) begin
                    if (4'h6 == idxUpdate_1[3:0]) begin
                      TBEMemory_6_way <= 3'h2;
                    end else begin
                      TBEMemory_6_way <= _GEN_455;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_6_way <= _GEN_455;
                    end else if (4'h6 == idxUpdate_1[3:0]) begin
                      TBEMemory_6_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_6_way <= _GEN_455;
                    end
                  end else begin
                    TBEMemory_6_way <= _GEN_455;
                  end
                end else if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEMemory_6_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_6_way <= _GEN_455;
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_way <= 3'h2;
                  end else begin
                    TBEMemory_6_way <= _GEN_455;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_6_way <= _GEN_455;
                  end else if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_6_way <= _GEN_455;
                  end
                end else begin
                  TBEMemory_6_way <= _GEN_455;
                end
              end else begin
                TBEMemory_6_way <= _GEN_969;
              end
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEMemory_6_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_6_way <= _GEN_969;
                end
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_way <= 3'h2;
                end else begin
                  TBEMemory_6_way <= _GEN_969;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_6_way <= _GEN_969;
                end else if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_6_way <= _GEN_969;
                end
              end else begin
                TBEMemory_6_way <= _GEN_969;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEMemory_6_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_6_way <= _GEN_969;
                  end
                end else if (_T_133) begin
                  if (4'h6 == idxUpdate_2[3:0]) begin
                    TBEMemory_6_way <= 3'h2;
                  end else begin
                    TBEMemory_6_way <= _GEN_969;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_6_way <= _GEN_969;
                  end else if (4'h6 == idxUpdate_2[3:0]) begin
                    TBEMemory_6_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_6_way <= _GEN_969;
                  end
                end else begin
                  TBEMemory_6_way <= _GEN_969;
                end
              end else if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEMemory_6_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_6_way <= _GEN_969;
                end
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_way <= 3'h2;
                end else begin
                  TBEMemory_6_way <= _GEN_969;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_6_way <= _GEN_969;
                end else if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_6_way <= _GEN_969;
                end
              end else begin
                TBEMemory_6_way <= _GEN_969;
              end
            end else begin
              TBEMemory_6_way <= _GEN_1483;
            end
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEMemory_6_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_6_way <= _GEN_1483;
              end
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_way <= 3'h2;
              end else begin
                TBEMemory_6_way <= _GEN_1483;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_6_way <= _GEN_1483;
              end else if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_6_way <= _GEN_1483;
              end
            end else begin
              TBEMemory_6_way <= _GEN_1483;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEMemory_6_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_6_way <= _GEN_1483;
                end
              end else if (_T_155) begin
                if (4'h6 == idxUpdate_3[3:0]) begin
                  TBEMemory_6_way <= 3'h2;
                end else begin
                  TBEMemory_6_way <= _GEN_1483;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_6_way <= _GEN_1483;
                end else if (4'h6 == idxUpdate_3[3:0]) begin
                  TBEMemory_6_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_6_way <= _GEN_1483;
                end
              end else begin
                TBEMemory_6_way <= _GEN_1483;
              end
            end else if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEMemory_6_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_6_way <= _GEN_1483;
              end
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_way <= 3'h2;
              end else begin
                TBEMemory_6_way <= _GEN_1483;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_6_way <= _GEN_1483;
              end else if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_6_way <= _GEN_1483;
              end
            end else begin
              TBEMemory_6_way <= _GEN_1483;
            end
          end else begin
            TBEMemory_6_way <= _GEN_1997;
          end
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEMemory_6_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_6_way <= _GEN_1997;
            end
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_way <= 3'h2;
            end else begin
              TBEMemory_6_way <= _GEN_1997;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_6_way <= _GEN_1997;
            end else if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_6_way <= _GEN_1997;
            end
          end else begin
            TBEMemory_6_way <= _GEN_1997;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEMemory_6_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_6_way <= _GEN_1997;
              end
            end else if (_T_177) begin
              if (4'h6 == idxUpdate_4[3:0]) begin
                TBEMemory_6_way <= 3'h2;
              end else begin
                TBEMemory_6_way <= _GEN_1997;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_6_way <= _GEN_1997;
              end else if (4'h6 == idxUpdate_4[3:0]) begin
                TBEMemory_6_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_6_way <= _GEN_1997;
              end
            end else begin
              TBEMemory_6_way <= _GEN_1997;
            end
          end else if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEMemory_6_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_6_way <= _GEN_1997;
            end
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_way <= 3'h2;
            end else begin
              TBEMemory_6_way <= _GEN_1997;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_6_way <= _GEN_1997;
            end else if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_6_way <= _GEN_1997;
            end
          end else begin
            TBEMemory_6_way <= _GEN_1997;
          end
        end else begin
          TBEMemory_6_way <= _GEN_2511;
        end
      end else if (_T_221) begin
        if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEMemory_6_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_6_way <= _GEN_2511;
          end
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_way <= 3'h2;
          end else begin
            TBEMemory_6_way <= _GEN_2511;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_6_way <= _GEN_2511;
          end else if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_6_way <= _GEN_2511;
          end
        end else begin
          TBEMemory_6_way <= _GEN_2511;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEMemory_6_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_6_way <= _GEN_2511;
            end
          end else if (_T_199) begin
            if (4'h6 == idxUpdate_5[3:0]) begin
              TBEMemory_6_way <= 3'h2;
            end else begin
              TBEMemory_6_way <= _GEN_2511;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_6_way <= _GEN_2511;
            end else if (4'h6 == idxUpdate_5[3:0]) begin
              TBEMemory_6_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_6_way <= _GEN_2511;
            end
          end else begin
            TBEMemory_6_way <= _GEN_2511;
          end
        end else if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEMemory_6_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_6_way <= _GEN_2511;
          end
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_way <= 3'h2;
          end else begin
            TBEMemory_6_way <= _GEN_2511;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_6_way <= _GEN_2511;
          end else if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_6_way <= _GEN_2511;
          end
        end else begin
          TBEMemory_6_way <= _GEN_2511;
        end
      end else begin
        TBEMemory_6_way <= _GEN_3025;
      end
    end else if (_T_243) begin
      if (4'h6 == idxUpdate_7[3:0]) begin
        TBEMemory_6_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'h6 == idxAlloc[3:0]) begin
          TBEMemory_6_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_6_way <= _GEN_3025;
        end
      end else if (_T_221) begin
        if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_way <= 3'h2;
        end else begin
          TBEMemory_6_way <= _GEN_3025;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_6_way <= _GEN_3025;
        end else if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_6_way <= _GEN_3025;
        end
      end else begin
        TBEMemory_6_way <= _GEN_3025;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEMemory_6_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_6_way <= _GEN_3025;
          end
        end else if (_T_221) begin
          if (4'h6 == idxUpdate_6[3:0]) begin
            TBEMemory_6_way <= 3'h2;
          end else begin
            TBEMemory_6_way <= _GEN_3025;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_6_way <= _GEN_3025;
          end else if (4'h6 == idxUpdate_6[3:0]) begin
            TBEMemory_6_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_6_way <= _GEN_3025;
          end
        end else begin
          TBEMemory_6_way <= _GEN_3025;
        end
      end else if (4'h6 == idxUpdate_7[3:0]) begin
        TBEMemory_6_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h6 == idxAlloc[3:0]) begin
          TBEMemory_6_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_6_way <= _GEN_3025;
        end
      end else if (_T_221) begin
        if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_way <= 3'h2;
        end else begin
          TBEMemory_6_way <= _GEN_3025;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_6_way <= _GEN_3025;
        end else if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_6_way <= _GEN_3025;
        end
      end else begin
        TBEMemory_6_way <= _GEN_3025;
      end
    end else begin
      TBEMemory_6_way <= _GEN_3539;
    end
    if (reset) begin
      TBEMemory_6_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h6 == idxAlloc[3:0]) begin
        TBEMemory_6_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'h6 == idxAlloc[3:0]) begin
          TBEMemory_6_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEMemory_6_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEMemory_6_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEMemory_6_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEMemory_6_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEMemory_6_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEMemory_6_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEMemory_6_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h6 == idxUpdate_0[3:0]) begin
                        TBEMemory_6_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEMemory_6_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEMemory_6_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h6 == idxUpdate_0[3:0]) begin
                        TBEMemory_6_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h6 == idxUpdate_1[3:0]) begin
                      TBEMemory_6_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'h6 == idxAlloc[3:0]) begin
                        TBEMemory_6_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'h6 == idxUpdate_0[3:0]) begin
                        TBEMemory_6_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'h6 == idxUpdate_0[3:0]) begin
                          TBEMemory_6_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEMemory_6_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEMemory_6_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h6 == idxUpdate_0[3:0]) begin
                        TBEMemory_6_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_439;
                end
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEMemory_6_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_439;
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_439;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h6 == idxUpdate_1[3:0]) begin
                      TBEMemory_6_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_6_fields_0 <= _GEN_439;
                    end
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_439;
                  end
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_439;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h6 == idxUpdate_2[3:0]) begin
                    TBEMemory_6_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEMemory_6_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_6_fields_0 <= _GEN_439;
                    end
                  end else if (_T_111) begin
                    if (4'h6 == idxUpdate_1[3:0]) begin
                      TBEMemory_6_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_6_fields_0 <= _GEN_439;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'h6 == idxUpdate_1[3:0]) begin
                        TBEMemory_6_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_6_fields_0 <= _GEN_439;
                      end
                    end else begin
                      TBEMemory_6_fields_0 <= _GEN_439;
                    end
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_439;
                  end
                end else if (isAlloc_1) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEMemory_6_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_439;
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEMemory_6_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_439;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h6 == idxUpdate_1[3:0]) begin
                      TBEMemory_6_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_6_fields_0 <= _GEN_439;
                    end
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_439;
                  end
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_439;
                end
              end else begin
                TBEMemory_6_fields_0 <= _GEN_953;
              end
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEMemory_6_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_953;
                end
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_953;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h6 == idxUpdate_2[3:0]) begin
                    TBEMemory_6_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_953;
                  end
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_953;
                end
              end else begin
                TBEMemory_6_fields_0 <= _GEN_953;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h6 == idxUpdate_3[3:0]) begin
                  TBEMemory_6_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEMemory_6_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_953;
                  end
                end else if (_T_133) begin
                  if (4'h6 == idxUpdate_2[3:0]) begin
                    TBEMemory_6_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_953;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'h6 == idxUpdate_2[3:0]) begin
                      TBEMemory_6_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_6_fields_0 <= _GEN_953;
                    end
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_953;
                  end
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_953;
                end
              end else if (isAlloc_2) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEMemory_6_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_953;
                end
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEMemory_6_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_953;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h6 == idxUpdate_2[3:0]) begin
                    TBEMemory_6_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_953;
                  end
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_953;
                end
              end else begin
                TBEMemory_6_fields_0 <= _GEN_953;
              end
            end else begin
              TBEMemory_6_fields_0 <= _GEN_1467;
            end
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEMemory_6_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_6_fields_0 <= _GEN_1467;
              end
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_fields_0 <= 32'h0;
              end else begin
                TBEMemory_6_fields_0 <= _GEN_1467;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h6 == idxUpdate_3[3:0]) begin
                  TBEMemory_6_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_1467;
                end
              end else begin
                TBEMemory_6_fields_0 <= _GEN_1467;
              end
            end else begin
              TBEMemory_6_fields_0 <= _GEN_1467;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h6 == idxUpdate_4[3:0]) begin
                TBEMemory_6_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEMemory_6_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_1467;
                end
              end else if (_T_155) begin
                if (4'h6 == idxUpdate_3[3:0]) begin
                  TBEMemory_6_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_1467;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'h6 == idxUpdate_3[3:0]) begin
                    TBEMemory_6_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_6_fields_0 <= _GEN_1467;
                  end
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_1467;
                end
              end else begin
                TBEMemory_6_fields_0 <= _GEN_1467;
              end
            end else if (isAlloc_3) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEMemory_6_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_6_fields_0 <= _GEN_1467;
              end
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEMemory_6_fields_0 <= 32'h0;
              end else begin
                TBEMemory_6_fields_0 <= _GEN_1467;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h6 == idxUpdate_3[3:0]) begin
                  TBEMemory_6_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_1467;
                end
              end else begin
                TBEMemory_6_fields_0 <= _GEN_1467;
              end
            end else begin
              TBEMemory_6_fields_0 <= _GEN_1467;
            end
          end else begin
            TBEMemory_6_fields_0 <= _GEN_1981;
          end
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEMemory_6_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_6_fields_0 <= _GEN_1981;
            end
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_fields_0 <= 32'h0;
            end else begin
              TBEMemory_6_fields_0 <= _GEN_1981;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h6 == idxUpdate_4[3:0]) begin
                TBEMemory_6_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_6_fields_0 <= _GEN_1981;
              end
            end else begin
              TBEMemory_6_fields_0 <= _GEN_1981;
            end
          end else begin
            TBEMemory_6_fields_0 <= _GEN_1981;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h6 == idxUpdate_5[3:0]) begin
              TBEMemory_6_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEMemory_6_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_6_fields_0 <= _GEN_1981;
              end
            end else if (_T_177) begin
              if (4'h6 == idxUpdate_4[3:0]) begin
                TBEMemory_6_fields_0 <= 32'h0;
              end else begin
                TBEMemory_6_fields_0 <= _GEN_1981;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'h6 == idxUpdate_4[3:0]) begin
                  TBEMemory_6_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_6_fields_0 <= _GEN_1981;
                end
              end else begin
                TBEMemory_6_fields_0 <= _GEN_1981;
              end
            end else begin
              TBEMemory_6_fields_0 <= _GEN_1981;
            end
          end else if (isAlloc_4) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEMemory_6_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_6_fields_0 <= _GEN_1981;
            end
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEMemory_6_fields_0 <= 32'h0;
            end else begin
              TBEMemory_6_fields_0 <= _GEN_1981;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h6 == idxUpdate_4[3:0]) begin
                TBEMemory_6_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_6_fields_0 <= _GEN_1981;
              end
            end else begin
              TBEMemory_6_fields_0 <= _GEN_1981;
            end
          end else begin
            TBEMemory_6_fields_0 <= _GEN_1981;
          end
        end else begin
          TBEMemory_6_fields_0 <= _GEN_2495;
        end
      end else if (_T_221) begin
        if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEMemory_6_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_6_fields_0 <= _GEN_2495;
          end
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_fields_0 <= 32'h0;
          end else begin
            TBEMemory_6_fields_0 <= _GEN_2495;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h6 == idxUpdate_5[3:0]) begin
              TBEMemory_6_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_6_fields_0 <= _GEN_2495;
            end
          end else begin
            TBEMemory_6_fields_0 <= _GEN_2495;
          end
        end else begin
          TBEMemory_6_fields_0 <= _GEN_2495;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h6 == idxUpdate_6[3:0]) begin
            TBEMemory_6_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEMemory_6_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_6_fields_0 <= _GEN_2495;
            end
          end else if (_T_199) begin
            if (4'h6 == idxUpdate_5[3:0]) begin
              TBEMemory_6_fields_0 <= 32'h0;
            end else begin
              TBEMemory_6_fields_0 <= _GEN_2495;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'h6 == idxUpdate_5[3:0]) begin
                TBEMemory_6_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_6_fields_0 <= _GEN_2495;
              end
            end else begin
              TBEMemory_6_fields_0 <= _GEN_2495;
            end
          end else begin
            TBEMemory_6_fields_0 <= _GEN_2495;
          end
        end else if (isAlloc_5) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEMemory_6_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_6_fields_0 <= _GEN_2495;
          end
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEMemory_6_fields_0 <= 32'h0;
          end else begin
            TBEMemory_6_fields_0 <= _GEN_2495;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h6 == idxUpdate_5[3:0]) begin
              TBEMemory_6_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_6_fields_0 <= _GEN_2495;
            end
          end else begin
            TBEMemory_6_fields_0 <= _GEN_2495;
          end
        end else begin
          TBEMemory_6_fields_0 <= _GEN_2495;
        end
      end else begin
        TBEMemory_6_fields_0 <= _GEN_3009;
      end
    end else if (_T_243) begin
      if (4'h6 == idxUpdate_7[3:0]) begin
        TBEMemory_6_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h6 == idxAlloc[3:0]) begin
          TBEMemory_6_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_6_fields_0 <= _GEN_3009;
        end
      end else if (_T_221) begin
        if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_fields_0 <= 32'h0;
        end else begin
          TBEMemory_6_fields_0 <= _GEN_3009;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h6 == idxUpdate_6[3:0]) begin
            TBEMemory_6_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_6_fields_0 <= _GEN_3009;
          end
        end else begin
          TBEMemory_6_fields_0 <= _GEN_3009;
        end
      end else begin
        TBEMemory_6_fields_0 <= _GEN_3009;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'h6 == idxUpdate_7[3:0]) begin
          TBEMemory_6_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEMemory_6_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_6_fields_0 <= _GEN_3009;
          end
        end else if (_T_221) begin
          if (4'h6 == idxUpdate_6[3:0]) begin
            TBEMemory_6_fields_0 <= 32'h0;
          end else begin
            TBEMemory_6_fields_0 <= _GEN_3009;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'h6 == idxUpdate_6[3:0]) begin
              TBEMemory_6_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_6_fields_0 <= _GEN_3009;
            end
          end else begin
            TBEMemory_6_fields_0 <= _GEN_3009;
          end
        end else begin
          TBEMemory_6_fields_0 <= _GEN_3009;
        end
      end else if (isAlloc_6) begin
        if (4'h6 == idxAlloc[3:0]) begin
          TBEMemory_6_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_6_fields_0 <= _GEN_3009;
        end
      end else if (_T_221) begin
        if (4'h6 == idxUpdate_6[3:0]) begin
          TBEMemory_6_fields_0 <= 32'h0;
        end else begin
          TBEMemory_6_fields_0 <= _GEN_3009;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h6 == idxUpdate_6[3:0]) begin
            TBEMemory_6_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_6_fields_0 <= _GEN_3009;
          end
        end else begin
          TBEMemory_6_fields_0 <= _GEN_3009;
        end
      end else begin
        TBEMemory_6_fields_0 <= _GEN_3009;
      end
    end else begin
      TBEMemory_6_fields_0 <= _GEN_3523;
    end
    if (reset) begin
      TBEMemory_7_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'h7 == idxAlloc[3:0]) begin
        TBEMemory_7_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h7 == idxAlloc[3:0]) begin
          TBEMemory_7_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEMemory_7_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEMemory_7_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEMemory_7_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEMemory_7_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEMemory_7_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEMemory_7_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEMemory_7_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h7 == idxUpdate_0[3:0]) begin
                        TBEMemory_7_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEMemory_7_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEMemory_7_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h7 == idxUpdate_0[3:0]) begin
                        TBEMemory_7_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h7 == idxAlloc[3:0]) begin
                        TBEMemory_7_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'h7 == idxUpdate_0[3:0]) begin
                        TBEMemory_7_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h7 == idxUpdate_0[3:0]) begin
                          TBEMemory_7_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEMemory_7_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEMemory_7_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h7 == idxUpdate_0[3:0]) begin
                        TBEMemory_7_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_7_state_state <= _GEN_472;
                end
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEMemory_7_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_7_state_state <= _GEN_472;
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_state_state <= 2'h0;
                  end else begin
                    TBEMemory_7_state_state <= _GEN_472;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_7_state_state <= _GEN_472;
                  end else if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_7_state_state <= _GEN_472;
                  end
                end else begin
                  TBEMemory_7_state_state <= _GEN_472;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEMemory_7_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_7_state_state <= _GEN_472;
                    end
                  end else if (_T_111) begin
                    if (4'h7 == idxUpdate_1[3:0]) begin
                      TBEMemory_7_state_state <= 2'h0;
                    end else begin
                      TBEMemory_7_state_state <= _GEN_472;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_7_state_state <= _GEN_472;
                    end else if (4'h7 == idxUpdate_1[3:0]) begin
                      TBEMemory_7_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_7_state_state <= _GEN_472;
                    end
                  end else begin
                    TBEMemory_7_state_state <= _GEN_472;
                  end
                end else if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEMemory_7_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_7_state_state <= _GEN_472;
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_state_state <= 2'h0;
                  end else begin
                    TBEMemory_7_state_state <= _GEN_472;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_7_state_state <= _GEN_472;
                  end else if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_7_state_state <= _GEN_472;
                  end
                end else begin
                  TBEMemory_7_state_state <= _GEN_472;
                end
              end else begin
                TBEMemory_7_state_state <= _GEN_986;
              end
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEMemory_7_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_7_state_state <= _GEN_986;
                end
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_state_state <= 2'h0;
                end else begin
                  TBEMemory_7_state_state <= _GEN_986;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_7_state_state <= _GEN_986;
                end else if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_7_state_state <= _GEN_986;
                end
              end else begin
                TBEMemory_7_state_state <= _GEN_986;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEMemory_7_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_7_state_state <= _GEN_986;
                  end
                end else if (_T_133) begin
                  if (4'h7 == idxUpdate_2[3:0]) begin
                    TBEMemory_7_state_state <= 2'h0;
                  end else begin
                    TBEMemory_7_state_state <= _GEN_986;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_7_state_state <= _GEN_986;
                  end else if (4'h7 == idxUpdate_2[3:0]) begin
                    TBEMemory_7_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_7_state_state <= _GEN_986;
                  end
                end else begin
                  TBEMemory_7_state_state <= _GEN_986;
                end
              end else if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEMemory_7_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_7_state_state <= _GEN_986;
                end
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_state_state <= 2'h0;
                end else begin
                  TBEMemory_7_state_state <= _GEN_986;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_7_state_state <= _GEN_986;
                end else if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_7_state_state <= _GEN_986;
                end
              end else begin
                TBEMemory_7_state_state <= _GEN_986;
              end
            end else begin
              TBEMemory_7_state_state <= _GEN_1500;
            end
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEMemory_7_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_7_state_state <= _GEN_1500;
              end
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_state_state <= 2'h0;
              end else begin
                TBEMemory_7_state_state <= _GEN_1500;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_7_state_state <= _GEN_1500;
              end else if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_7_state_state <= _GEN_1500;
              end
            end else begin
              TBEMemory_7_state_state <= _GEN_1500;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEMemory_7_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_7_state_state <= _GEN_1500;
                end
              end else if (_T_155) begin
                if (4'h7 == idxUpdate_3[3:0]) begin
                  TBEMemory_7_state_state <= 2'h0;
                end else begin
                  TBEMemory_7_state_state <= _GEN_1500;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_7_state_state <= _GEN_1500;
                end else if (4'h7 == idxUpdate_3[3:0]) begin
                  TBEMemory_7_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_7_state_state <= _GEN_1500;
                end
              end else begin
                TBEMemory_7_state_state <= _GEN_1500;
              end
            end else if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEMemory_7_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_7_state_state <= _GEN_1500;
              end
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_state_state <= 2'h0;
              end else begin
                TBEMemory_7_state_state <= _GEN_1500;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_7_state_state <= _GEN_1500;
              end else if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_7_state_state <= _GEN_1500;
              end
            end else begin
              TBEMemory_7_state_state <= _GEN_1500;
            end
          end else begin
            TBEMemory_7_state_state <= _GEN_2014;
          end
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEMemory_7_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_7_state_state <= _GEN_2014;
            end
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_state_state <= 2'h0;
            end else begin
              TBEMemory_7_state_state <= _GEN_2014;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_7_state_state <= _GEN_2014;
            end else if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_7_state_state <= _GEN_2014;
            end
          end else begin
            TBEMemory_7_state_state <= _GEN_2014;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEMemory_7_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_7_state_state <= _GEN_2014;
              end
            end else if (_T_177) begin
              if (4'h7 == idxUpdate_4[3:0]) begin
                TBEMemory_7_state_state <= 2'h0;
              end else begin
                TBEMemory_7_state_state <= _GEN_2014;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_7_state_state <= _GEN_2014;
              end else if (4'h7 == idxUpdate_4[3:0]) begin
                TBEMemory_7_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_7_state_state <= _GEN_2014;
              end
            end else begin
              TBEMemory_7_state_state <= _GEN_2014;
            end
          end else if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEMemory_7_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_7_state_state <= _GEN_2014;
            end
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_state_state <= 2'h0;
            end else begin
              TBEMemory_7_state_state <= _GEN_2014;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_7_state_state <= _GEN_2014;
            end else if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_7_state_state <= _GEN_2014;
            end
          end else begin
            TBEMemory_7_state_state <= _GEN_2014;
          end
        end else begin
          TBEMemory_7_state_state <= _GEN_2528;
        end
      end else if (_T_221) begin
        if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEMemory_7_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_7_state_state <= _GEN_2528;
          end
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_state_state <= 2'h0;
          end else begin
            TBEMemory_7_state_state <= _GEN_2528;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_7_state_state <= _GEN_2528;
          end else if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_7_state_state <= _GEN_2528;
          end
        end else begin
          TBEMemory_7_state_state <= _GEN_2528;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEMemory_7_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_7_state_state <= _GEN_2528;
            end
          end else if (_T_199) begin
            if (4'h7 == idxUpdate_5[3:0]) begin
              TBEMemory_7_state_state <= 2'h0;
            end else begin
              TBEMemory_7_state_state <= _GEN_2528;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_7_state_state <= _GEN_2528;
            end else if (4'h7 == idxUpdate_5[3:0]) begin
              TBEMemory_7_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_7_state_state <= _GEN_2528;
            end
          end else begin
            TBEMemory_7_state_state <= _GEN_2528;
          end
        end else if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEMemory_7_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_7_state_state <= _GEN_2528;
          end
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_state_state <= 2'h0;
          end else begin
            TBEMemory_7_state_state <= _GEN_2528;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_7_state_state <= _GEN_2528;
          end else if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_7_state_state <= _GEN_2528;
          end
        end else begin
          TBEMemory_7_state_state <= _GEN_2528;
        end
      end else begin
        TBEMemory_7_state_state <= _GEN_3042;
      end
    end else if (_T_243) begin
      if (4'h7 == idxUpdate_7[3:0]) begin
        TBEMemory_7_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'h7 == idxAlloc[3:0]) begin
          TBEMemory_7_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_7_state_state <= _GEN_3042;
        end
      end else if (_T_221) begin
        if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_state_state <= 2'h0;
        end else begin
          TBEMemory_7_state_state <= _GEN_3042;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_7_state_state <= _GEN_3042;
        end else if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_7_state_state <= _GEN_3042;
        end
      end else begin
        TBEMemory_7_state_state <= _GEN_3042;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEMemory_7_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_7_state_state <= _GEN_3042;
          end
        end else if (_T_221) begin
          if (4'h7 == idxUpdate_6[3:0]) begin
            TBEMemory_7_state_state <= 2'h0;
          end else begin
            TBEMemory_7_state_state <= _GEN_3042;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_7_state_state <= _GEN_3042;
          end else if (4'h7 == idxUpdate_6[3:0]) begin
            TBEMemory_7_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_7_state_state <= _GEN_3042;
          end
        end else begin
          TBEMemory_7_state_state <= _GEN_3042;
        end
      end else if (4'h7 == idxUpdate_7[3:0]) begin
        TBEMemory_7_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h7 == idxAlloc[3:0]) begin
          TBEMemory_7_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_7_state_state <= _GEN_3042;
        end
      end else if (_T_221) begin
        if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_state_state <= 2'h0;
        end else begin
          TBEMemory_7_state_state <= _GEN_3042;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_7_state_state <= _GEN_3042;
        end else if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_7_state_state <= _GEN_3042;
        end
      end else begin
        TBEMemory_7_state_state <= _GEN_3042;
      end
    end else begin
      TBEMemory_7_state_state <= _GEN_3556;
    end
    if (reset) begin
      TBEMemory_7_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'h7 == idxAlloc[3:0]) begin
        TBEMemory_7_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h7 == idxAlloc[3:0]) begin
          TBEMemory_7_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEMemory_7_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEMemory_7_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEMemory_7_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEMemory_7_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEMemory_7_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEMemory_7_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEMemory_7_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h7 == idxUpdate_0[3:0]) begin
                        TBEMemory_7_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEMemory_7_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEMemory_7_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h7 == idxUpdate_0[3:0]) begin
                        TBEMemory_7_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h7 == idxAlloc[3:0]) begin
                        TBEMemory_7_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'h7 == idxUpdate_0[3:0]) begin
                        TBEMemory_7_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h7 == idxUpdate_0[3:0]) begin
                          TBEMemory_7_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEMemory_7_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEMemory_7_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h7 == idxUpdate_0[3:0]) begin
                        TBEMemory_7_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_7_way <= _GEN_456;
                end
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEMemory_7_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_7_way <= _GEN_456;
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_way <= 3'h2;
                  end else begin
                    TBEMemory_7_way <= _GEN_456;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_7_way <= _GEN_456;
                  end else if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_7_way <= _GEN_456;
                  end
                end else begin
                  TBEMemory_7_way <= _GEN_456;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEMemory_7_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_7_way <= _GEN_456;
                    end
                  end else if (_T_111) begin
                    if (4'h7 == idxUpdate_1[3:0]) begin
                      TBEMemory_7_way <= 3'h2;
                    end else begin
                      TBEMemory_7_way <= _GEN_456;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_7_way <= _GEN_456;
                    end else if (4'h7 == idxUpdate_1[3:0]) begin
                      TBEMemory_7_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_7_way <= _GEN_456;
                    end
                  end else begin
                    TBEMemory_7_way <= _GEN_456;
                  end
                end else if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEMemory_7_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_7_way <= _GEN_456;
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_way <= 3'h2;
                  end else begin
                    TBEMemory_7_way <= _GEN_456;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_7_way <= _GEN_456;
                  end else if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_7_way <= _GEN_456;
                  end
                end else begin
                  TBEMemory_7_way <= _GEN_456;
                end
              end else begin
                TBEMemory_7_way <= _GEN_970;
              end
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEMemory_7_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_7_way <= _GEN_970;
                end
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_way <= 3'h2;
                end else begin
                  TBEMemory_7_way <= _GEN_970;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_7_way <= _GEN_970;
                end else if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_7_way <= _GEN_970;
                end
              end else begin
                TBEMemory_7_way <= _GEN_970;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEMemory_7_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_7_way <= _GEN_970;
                  end
                end else if (_T_133) begin
                  if (4'h7 == idxUpdate_2[3:0]) begin
                    TBEMemory_7_way <= 3'h2;
                  end else begin
                    TBEMemory_7_way <= _GEN_970;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_7_way <= _GEN_970;
                  end else if (4'h7 == idxUpdate_2[3:0]) begin
                    TBEMemory_7_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_7_way <= _GEN_970;
                  end
                end else begin
                  TBEMemory_7_way <= _GEN_970;
                end
              end else if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEMemory_7_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_7_way <= _GEN_970;
                end
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_way <= 3'h2;
                end else begin
                  TBEMemory_7_way <= _GEN_970;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_7_way <= _GEN_970;
                end else if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_7_way <= _GEN_970;
                end
              end else begin
                TBEMemory_7_way <= _GEN_970;
              end
            end else begin
              TBEMemory_7_way <= _GEN_1484;
            end
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEMemory_7_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_7_way <= _GEN_1484;
              end
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_way <= 3'h2;
              end else begin
                TBEMemory_7_way <= _GEN_1484;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_7_way <= _GEN_1484;
              end else if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_7_way <= _GEN_1484;
              end
            end else begin
              TBEMemory_7_way <= _GEN_1484;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEMemory_7_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_7_way <= _GEN_1484;
                end
              end else if (_T_155) begin
                if (4'h7 == idxUpdate_3[3:0]) begin
                  TBEMemory_7_way <= 3'h2;
                end else begin
                  TBEMemory_7_way <= _GEN_1484;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_7_way <= _GEN_1484;
                end else if (4'h7 == idxUpdate_3[3:0]) begin
                  TBEMemory_7_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_7_way <= _GEN_1484;
                end
              end else begin
                TBEMemory_7_way <= _GEN_1484;
              end
            end else if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEMemory_7_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_7_way <= _GEN_1484;
              end
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_way <= 3'h2;
              end else begin
                TBEMemory_7_way <= _GEN_1484;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_7_way <= _GEN_1484;
              end else if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_7_way <= _GEN_1484;
              end
            end else begin
              TBEMemory_7_way <= _GEN_1484;
            end
          end else begin
            TBEMemory_7_way <= _GEN_1998;
          end
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEMemory_7_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_7_way <= _GEN_1998;
            end
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_way <= 3'h2;
            end else begin
              TBEMemory_7_way <= _GEN_1998;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_7_way <= _GEN_1998;
            end else if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_7_way <= _GEN_1998;
            end
          end else begin
            TBEMemory_7_way <= _GEN_1998;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEMemory_7_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_7_way <= _GEN_1998;
              end
            end else if (_T_177) begin
              if (4'h7 == idxUpdate_4[3:0]) begin
                TBEMemory_7_way <= 3'h2;
              end else begin
                TBEMemory_7_way <= _GEN_1998;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_7_way <= _GEN_1998;
              end else if (4'h7 == idxUpdate_4[3:0]) begin
                TBEMemory_7_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_7_way <= _GEN_1998;
              end
            end else begin
              TBEMemory_7_way <= _GEN_1998;
            end
          end else if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEMemory_7_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_7_way <= _GEN_1998;
            end
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_way <= 3'h2;
            end else begin
              TBEMemory_7_way <= _GEN_1998;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_7_way <= _GEN_1998;
            end else if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_7_way <= _GEN_1998;
            end
          end else begin
            TBEMemory_7_way <= _GEN_1998;
          end
        end else begin
          TBEMemory_7_way <= _GEN_2512;
        end
      end else if (_T_221) begin
        if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEMemory_7_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_7_way <= _GEN_2512;
          end
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_way <= 3'h2;
          end else begin
            TBEMemory_7_way <= _GEN_2512;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_7_way <= _GEN_2512;
          end else if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_7_way <= _GEN_2512;
          end
        end else begin
          TBEMemory_7_way <= _GEN_2512;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEMemory_7_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_7_way <= _GEN_2512;
            end
          end else if (_T_199) begin
            if (4'h7 == idxUpdate_5[3:0]) begin
              TBEMemory_7_way <= 3'h2;
            end else begin
              TBEMemory_7_way <= _GEN_2512;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_7_way <= _GEN_2512;
            end else if (4'h7 == idxUpdate_5[3:0]) begin
              TBEMemory_7_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_7_way <= _GEN_2512;
            end
          end else begin
            TBEMemory_7_way <= _GEN_2512;
          end
        end else if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEMemory_7_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_7_way <= _GEN_2512;
          end
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_way <= 3'h2;
          end else begin
            TBEMemory_7_way <= _GEN_2512;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_7_way <= _GEN_2512;
          end else if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_7_way <= _GEN_2512;
          end
        end else begin
          TBEMemory_7_way <= _GEN_2512;
        end
      end else begin
        TBEMemory_7_way <= _GEN_3026;
      end
    end else if (_T_243) begin
      if (4'h7 == idxUpdate_7[3:0]) begin
        TBEMemory_7_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'h7 == idxAlloc[3:0]) begin
          TBEMemory_7_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_7_way <= _GEN_3026;
        end
      end else if (_T_221) begin
        if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_way <= 3'h2;
        end else begin
          TBEMemory_7_way <= _GEN_3026;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_7_way <= _GEN_3026;
        end else if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_7_way <= _GEN_3026;
        end
      end else begin
        TBEMemory_7_way <= _GEN_3026;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEMemory_7_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_7_way <= _GEN_3026;
          end
        end else if (_T_221) begin
          if (4'h7 == idxUpdate_6[3:0]) begin
            TBEMemory_7_way <= 3'h2;
          end else begin
            TBEMemory_7_way <= _GEN_3026;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_7_way <= _GEN_3026;
          end else if (4'h7 == idxUpdate_6[3:0]) begin
            TBEMemory_7_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_7_way <= _GEN_3026;
          end
        end else begin
          TBEMemory_7_way <= _GEN_3026;
        end
      end else if (4'h7 == idxUpdate_7[3:0]) begin
        TBEMemory_7_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h7 == idxAlloc[3:0]) begin
          TBEMemory_7_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_7_way <= _GEN_3026;
        end
      end else if (_T_221) begin
        if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_way <= 3'h2;
        end else begin
          TBEMemory_7_way <= _GEN_3026;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_7_way <= _GEN_3026;
        end else if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_7_way <= _GEN_3026;
        end
      end else begin
        TBEMemory_7_way <= _GEN_3026;
      end
    end else begin
      TBEMemory_7_way <= _GEN_3540;
    end
    if (reset) begin
      TBEMemory_7_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h7 == idxAlloc[3:0]) begin
        TBEMemory_7_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'h7 == idxAlloc[3:0]) begin
          TBEMemory_7_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEMemory_7_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEMemory_7_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEMemory_7_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEMemory_7_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEMemory_7_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEMemory_7_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEMemory_7_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h7 == idxUpdate_0[3:0]) begin
                        TBEMemory_7_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEMemory_7_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEMemory_7_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h7 == idxUpdate_0[3:0]) begin
                        TBEMemory_7_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h7 == idxUpdate_1[3:0]) begin
                      TBEMemory_7_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'h7 == idxAlloc[3:0]) begin
                        TBEMemory_7_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'h7 == idxUpdate_0[3:0]) begin
                        TBEMemory_7_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'h7 == idxUpdate_0[3:0]) begin
                          TBEMemory_7_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEMemory_7_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEMemory_7_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h7 == idxUpdate_0[3:0]) begin
                        TBEMemory_7_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_440;
                end
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEMemory_7_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_440;
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_440;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h7 == idxUpdate_1[3:0]) begin
                      TBEMemory_7_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_7_fields_0 <= _GEN_440;
                    end
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_440;
                  end
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_440;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h7 == idxUpdate_2[3:0]) begin
                    TBEMemory_7_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEMemory_7_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_7_fields_0 <= _GEN_440;
                    end
                  end else if (_T_111) begin
                    if (4'h7 == idxUpdate_1[3:0]) begin
                      TBEMemory_7_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_7_fields_0 <= _GEN_440;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'h7 == idxUpdate_1[3:0]) begin
                        TBEMemory_7_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_7_fields_0 <= _GEN_440;
                      end
                    end else begin
                      TBEMemory_7_fields_0 <= _GEN_440;
                    end
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_440;
                  end
                end else if (isAlloc_1) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEMemory_7_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_440;
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEMemory_7_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_440;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h7 == idxUpdate_1[3:0]) begin
                      TBEMemory_7_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_7_fields_0 <= _GEN_440;
                    end
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_440;
                  end
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_440;
                end
              end else begin
                TBEMemory_7_fields_0 <= _GEN_954;
              end
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEMemory_7_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_954;
                end
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_954;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h7 == idxUpdate_2[3:0]) begin
                    TBEMemory_7_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_954;
                  end
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_954;
                end
              end else begin
                TBEMemory_7_fields_0 <= _GEN_954;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h7 == idxUpdate_3[3:0]) begin
                  TBEMemory_7_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEMemory_7_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_954;
                  end
                end else if (_T_133) begin
                  if (4'h7 == idxUpdate_2[3:0]) begin
                    TBEMemory_7_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_954;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'h7 == idxUpdate_2[3:0]) begin
                      TBEMemory_7_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_7_fields_0 <= _GEN_954;
                    end
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_954;
                  end
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_954;
                end
              end else if (isAlloc_2) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEMemory_7_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_954;
                end
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEMemory_7_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_954;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h7 == idxUpdate_2[3:0]) begin
                    TBEMemory_7_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_954;
                  end
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_954;
                end
              end else begin
                TBEMemory_7_fields_0 <= _GEN_954;
              end
            end else begin
              TBEMemory_7_fields_0 <= _GEN_1468;
            end
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEMemory_7_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_7_fields_0 <= _GEN_1468;
              end
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_fields_0 <= 32'h0;
              end else begin
                TBEMemory_7_fields_0 <= _GEN_1468;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h7 == idxUpdate_3[3:0]) begin
                  TBEMemory_7_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_1468;
                end
              end else begin
                TBEMemory_7_fields_0 <= _GEN_1468;
              end
            end else begin
              TBEMemory_7_fields_0 <= _GEN_1468;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h7 == idxUpdate_4[3:0]) begin
                TBEMemory_7_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEMemory_7_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_1468;
                end
              end else if (_T_155) begin
                if (4'h7 == idxUpdate_3[3:0]) begin
                  TBEMemory_7_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_1468;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'h7 == idxUpdate_3[3:0]) begin
                    TBEMemory_7_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_7_fields_0 <= _GEN_1468;
                  end
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_1468;
                end
              end else begin
                TBEMemory_7_fields_0 <= _GEN_1468;
              end
            end else if (isAlloc_3) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEMemory_7_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_7_fields_0 <= _GEN_1468;
              end
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEMemory_7_fields_0 <= 32'h0;
              end else begin
                TBEMemory_7_fields_0 <= _GEN_1468;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h7 == idxUpdate_3[3:0]) begin
                  TBEMemory_7_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_1468;
                end
              end else begin
                TBEMemory_7_fields_0 <= _GEN_1468;
              end
            end else begin
              TBEMemory_7_fields_0 <= _GEN_1468;
            end
          end else begin
            TBEMemory_7_fields_0 <= _GEN_1982;
          end
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEMemory_7_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_7_fields_0 <= _GEN_1982;
            end
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_fields_0 <= 32'h0;
            end else begin
              TBEMemory_7_fields_0 <= _GEN_1982;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h7 == idxUpdate_4[3:0]) begin
                TBEMemory_7_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_7_fields_0 <= _GEN_1982;
              end
            end else begin
              TBEMemory_7_fields_0 <= _GEN_1982;
            end
          end else begin
            TBEMemory_7_fields_0 <= _GEN_1982;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h7 == idxUpdate_5[3:0]) begin
              TBEMemory_7_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEMemory_7_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_7_fields_0 <= _GEN_1982;
              end
            end else if (_T_177) begin
              if (4'h7 == idxUpdate_4[3:0]) begin
                TBEMemory_7_fields_0 <= 32'h0;
              end else begin
                TBEMemory_7_fields_0 <= _GEN_1982;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'h7 == idxUpdate_4[3:0]) begin
                  TBEMemory_7_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_7_fields_0 <= _GEN_1982;
                end
              end else begin
                TBEMemory_7_fields_0 <= _GEN_1982;
              end
            end else begin
              TBEMemory_7_fields_0 <= _GEN_1982;
            end
          end else if (isAlloc_4) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEMemory_7_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_7_fields_0 <= _GEN_1982;
            end
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEMemory_7_fields_0 <= 32'h0;
            end else begin
              TBEMemory_7_fields_0 <= _GEN_1982;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h7 == idxUpdate_4[3:0]) begin
                TBEMemory_7_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_7_fields_0 <= _GEN_1982;
              end
            end else begin
              TBEMemory_7_fields_0 <= _GEN_1982;
            end
          end else begin
            TBEMemory_7_fields_0 <= _GEN_1982;
          end
        end else begin
          TBEMemory_7_fields_0 <= _GEN_2496;
        end
      end else if (_T_221) begin
        if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEMemory_7_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_7_fields_0 <= _GEN_2496;
          end
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_fields_0 <= 32'h0;
          end else begin
            TBEMemory_7_fields_0 <= _GEN_2496;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h7 == idxUpdate_5[3:0]) begin
              TBEMemory_7_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_7_fields_0 <= _GEN_2496;
            end
          end else begin
            TBEMemory_7_fields_0 <= _GEN_2496;
          end
        end else begin
          TBEMemory_7_fields_0 <= _GEN_2496;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h7 == idxUpdate_6[3:0]) begin
            TBEMemory_7_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEMemory_7_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_7_fields_0 <= _GEN_2496;
            end
          end else if (_T_199) begin
            if (4'h7 == idxUpdate_5[3:0]) begin
              TBEMemory_7_fields_0 <= 32'h0;
            end else begin
              TBEMemory_7_fields_0 <= _GEN_2496;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'h7 == idxUpdate_5[3:0]) begin
                TBEMemory_7_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_7_fields_0 <= _GEN_2496;
              end
            end else begin
              TBEMemory_7_fields_0 <= _GEN_2496;
            end
          end else begin
            TBEMemory_7_fields_0 <= _GEN_2496;
          end
        end else if (isAlloc_5) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEMemory_7_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_7_fields_0 <= _GEN_2496;
          end
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEMemory_7_fields_0 <= 32'h0;
          end else begin
            TBEMemory_7_fields_0 <= _GEN_2496;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h7 == idxUpdate_5[3:0]) begin
              TBEMemory_7_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_7_fields_0 <= _GEN_2496;
            end
          end else begin
            TBEMemory_7_fields_0 <= _GEN_2496;
          end
        end else begin
          TBEMemory_7_fields_0 <= _GEN_2496;
        end
      end else begin
        TBEMemory_7_fields_0 <= _GEN_3010;
      end
    end else if (_T_243) begin
      if (4'h7 == idxUpdate_7[3:0]) begin
        TBEMemory_7_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h7 == idxAlloc[3:0]) begin
          TBEMemory_7_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_7_fields_0 <= _GEN_3010;
        end
      end else if (_T_221) begin
        if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_fields_0 <= 32'h0;
        end else begin
          TBEMemory_7_fields_0 <= _GEN_3010;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h7 == idxUpdate_6[3:0]) begin
            TBEMemory_7_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_7_fields_0 <= _GEN_3010;
          end
        end else begin
          TBEMemory_7_fields_0 <= _GEN_3010;
        end
      end else begin
        TBEMemory_7_fields_0 <= _GEN_3010;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'h7 == idxUpdate_7[3:0]) begin
          TBEMemory_7_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEMemory_7_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_7_fields_0 <= _GEN_3010;
          end
        end else if (_T_221) begin
          if (4'h7 == idxUpdate_6[3:0]) begin
            TBEMemory_7_fields_0 <= 32'h0;
          end else begin
            TBEMemory_7_fields_0 <= _GEN_3010;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'h7 == idxUpdate_6[3:0]) begin
              TBEMemory_7_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_7_fields_0 <= _GEN_3010;
            end
          end else begin
            TBEMemory_7_fields_0 <= _GEN_3010;
          end
        end else begin
          TBEMemory_7_fields_0 <= _GEN_3010;
        end
      end else if (isAlloc_6) begin
        if (4'h7 == idxAlloc[3:0]) begin
          TBEMemory_7_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_7_fields_0 <= _GEN_3010;
        end
      end else if (_T_221) begin
        if (4'h7 == idxUpdate_6[3:0]) begin
          TBEMemory_7_fields_0 <= 32'h0;
        end else begin
          TBEMemory_7_fields_0 <= _GEN_3010;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h7 == idxUpdate_6[3:0]) begin
            TBEMemory_7_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_7_fields_0 <= _GEN_3010;
          end
        end else begin
          TBEMemory_7_fields_0 <= _GEN_3010;
        end
      end else begin
        TBEMemory_7_fields_0 <= _GEN_3010;
      end
    end else begin
      TBEMemory_7_fields_0 <= _GEN_3524;
    end
    if (reset) begin
      TBEMemory_8_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'h8 == idxAlloc[3:0]) begin
        TBEMemory_8_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h8 == idxAlloc[3:0]) begin
          TBEMemory_8_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEMemory_8_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEMemory_8_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEMemory_8_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEMemory_8_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEMemory_8_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEMemory_8_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEMemory_8_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h8 == idxUpdate_0[3:0]) begin
                        TBEMemory_8_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEMemory_8_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEMemory_8_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h8 == idxUpdate_0[3:0]) begin
                        TBEMemory_8_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h8 == idxAlloc[3:0]) begin
                        TBEMemory_8_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'h8 == idxUpdate_0[3:0]) begin
                        TBEMemory_8_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h8 == idxUpdate_0[3:0]) begin
                          TBEMemory_8_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEMemory_8_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEMemory_8_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h8 == idxUpdate_0[3:0]) begin
                        TBEMemory_8_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_8_state_state <= _GEN_473;
                end
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEMemory_8_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_8_state_state <= _GEN_473;
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_state_state <= 2'h0;
                  end else begin
                    TBEMemory_8_state_state <= _GEN_473;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_8_state_state <= _GEN_473;
                  end else if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_8_state_state <= _GEN_473;
                  end
                end else begin
                  TBEMemory_8_state_state <= _GEN_473;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEMemory_8_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_8_state_state <= _GEN_473;
                    end
                  end else if (_T_111) begin
                    if (4'h8 == idxUpdate_1[3:0]) begin
                      TBEMemory_8_state_state <= 2'h0;
                    end else begin
                      TBEMemory_8_state_state <= _GEN_473;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_8_state_state <= _GEN_473;
                    end else if (4'h8 == idxUpdate_1[3:0]) begin
                      TBEMemory_8_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_8_state_state <= _GEN_473;
                    end
                  end else begin
                    TBEMemory_8_state_state <= _GEN_473;
                  end
                end else if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEMemory_8_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_8_state_state <= _GEN_473;
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_state_state <= 2'h0;
                  end else begin
                    TBEMemory_8_state_state <= _GEN_473;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_8_state_state <= _GEN_473;
                  end else if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_8_state_state <= _GEN_473;
                  end
                end else begin
                  TBEMemory_8_state_state <= _GEN_473;
                end
              end else begin
                TBEMemory_8_state_state <= _GEN_987;
              end
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEMemory_8_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_8_state_state <= _GEN_987;
                end
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_state_state <= 2'h0;
                end else begin
                  TBEMemory_8_state_state <= _GEN_987;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_8_state_state <= _GEN_987;
                end else if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_8_state_state <= _GEN_987;
                end
              end else begin
                TBEMemory_8_state_state <= _GEN_987;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEMemory_8_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_8_state_state <= _GEN_987;
                  end
                end else if (_T_133) begin
                  if (4'h8 == idxUpdate_2[3:0]) begin
                    TBEMemory_8_state_state <= 2'h0;
                  end else begin
                    TBEMemory_8_state_state <= _GEN_987;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_8_state_state <= _GEN_987;
                  end else if (4'h8 == idxUpdate_2[3:0]) begin
                    TBEMemory_8_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_8_state_state <= _GEN_987;
                  end
                end else begin
                  TBEMemory_8_state_state <= _GEN_987;
                end
              end else if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEMemory_8_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_8_state_state <= _GEN_987;
                end
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_state_state <= 2'h0;
                end else begin
                  TBEMemory_8_state_state <= _GEN_987;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_8_state_state <= _GEN_987;
                end else if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_8_state_state <= _GEN_987;
                end
              end else begin
                TBEMemory_8_state_state <= _GEN_987;
              end
            end else begin
              TBEMemory_8_state_state <= _GEN_1501;
            end
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEMemory_8_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_8_state_state <= _GEN_1501;
              end
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_state_state <= 2'h0;
              end else begin
                TBEMemory_8_state_state <= _GEN_1501;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_8_state_state <= _GEN_1501;
              end else if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_8_state_state <= _GEN_1501;
              end
            end else begin
              TBEMemory_8_state_state <= _GEN_1501;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEMemory_8_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_8_state_state <= _GEN_1501;
                end
              end else if (_T_155) begin
                if (4'h8 == idxUpdate_3[3:0]) begin
                  TBEMemory_8_state_state <= 2'h0;
                end else begin
                  TBEMemory_8_state_state <= _GEN_1501;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_8_state_state <= _GEN_1501;
                end else if (4'h8 == idxUpdate_3[3:0]) begin
                  TBEMemory_8_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_8_state_state <= _GEN_1501;
                end
              end else begin
                TBEMemory_8_state_state <= _GEN_1501;
              end
            end else if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEMemory_8_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_8_state_state <= _GEN_1501;
              end
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_state_state <= 2'h0;
              end else begin
                TBEMemory_8_state_state <= _GEN_1501;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_8_state_state <= _GEN_1501;
              end else if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_8_state_state <= _GEN_1501;
              end
            end else begin
              TBEMemory_8_state_state <= _GEN_1501;
            end
          end else begin
            TBEMemory_8_state_state <= _GEN_2015;
          end
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEMemory_8_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_8_state_state <= _GEN_2015;
            end
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_state_state <= 2'h0;
            end else begin
              TBEMemory_8_state_state <= _GEN_2015;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_8_state_state <= _GEN_2015;
            end else if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_8_state_state <= _GEN_2015;
            end
          end else begin
            TBEMemory_8_state_state <= _GEN_2015;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEMemory_8_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_8_state_state <= _GEN_2015;
              end
            end else if (_T_177) begin
              if (4'h8 == idxUpdate_4[3:0]) begin
                TBEMemory_8_state_state <= 2'h0;
              end else begin
                TBEMemory_8_state_state <= _GEN_2015;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_8_state_state <= _GEN_2015;
              end else if (4'h8 == idxUpdate_4[3:0]) begin
                TBEMemory_8_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_8_state_state <= _GEN_2015;
              end
            end else begin
              TBEMemory_8_state_state <= _GEN_2015;
            end
          end else if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEMemory_8_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_8_state_state <= _GEN_2015;
            end
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_state_state <= 2'h0;
            end else begin
              TBEMemory_8_state_state <= _GEN_2015;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_8_state_state <= _GEN_2015;
            end else if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_8_state_state <= _GEN_2015;
            end
          end else begin
            TBEMemory_8_state_state <= _GEN_2015;
          end
        end else begin
          TBEMemory_8_state_state <= _GEN_2529;
        end
      end else if (_T_221) begin
        if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEMemory_8_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_8_state_state <= _GEN_2529;
          end
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_state_state <= 2'h0;
          end else begin
            TBEMemory_8_state_state <= _GEN_2529;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_8_state_state <= _GEN_2529;
          end else if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_8_state_state <= _GEN_2529;
          end
        end else begin
          TBEMemory_8_state_state <= _GEN_2529;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEMemory_8_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_8_state_state <= _GEN_2529;
            end
          end else if (_T_199) begin
            if (4'h8 == idxUpdate_5[3:0]) begin
              TBEMemory_8_state_state <= 2'h0;
            end else begin
              TBEMemory_8_state_state <= _GEN_2529;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_8_state_state <= _GEN_2529;
            end else if (4'h8 == idxUpdate_5[3:0]) begin
              TBEMemory_8_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_8_state_state <= _GEN_2529;
            end
          end else begin
            TBEMemory_8_state_state <= _GEN_2529;
          end
        end else if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEMemory_8_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_8_state_state <= _GEN_2529;
          end
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_state_state <= 2'h0;
          end else begin
            TBEMemory_8_state_state <= _GEN_2529;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_8_state_state <= _GEN_2529;
          end else if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_8_state_state <= _GEN_2529;
          end
        end else begin
          TBEMemory_8_state_state <= _GEN_2529;
        end
      end else begin
        TBEMemory_8_state_state <= _GEN_3043;
      end
    end else if (_T_243) begin
      if (4'h8 == idxUpdate_7[3:0]) begin
        TBEMemory_8_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'h8 == idxAlloc[3:0]) begin
          TBEMemory_8_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_8_state_state <= _GEN_3043;
        end
      end else if (_T_221) begin
        if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_state_state <= 2'h0;
        end else begin
          TBEMemory_8_state_state <= _GEN_3043;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_8_state_state <= _GEN_3043;
        end else if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_8_state_state <= _GEN_3043;
        end
      end else begin
        TBEMemory_8_state_state <= _GEN_3043;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEMemory_8_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_8_state_state <= _GEN_3043;
          end
        end else if (_T_221) begin
          if (4'h8 == idxUpdate_6[3:0]) begin
            TBEMemory_8_state_state <= 2'h0;
          end else begin
            TBEMemory_8_state_state <= _GEN_3043;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_8_state_state <= _GEN_3043;
          end else if (4'h8 == idxUpdate_6[3:0]) begin
            TBEMemory_8_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_8_state_state <= _GEN_3043;
          end
        end else begin
          TBEMemory_8_state_state <= _GEN_3043;
        end
      end else if (4'h8 == idxUpdate_7[3:0]) begin
        TBEMemory_8_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h8 == idxAlloc[3:0]) begin
          TBEMemory_8_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_8_state_state <= _GEN_3043;
        end
      end else if (_T_221) begin
        if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_state_state <= 2'h0;
        end else begin
          TBEMemory_8_state_state <= _GEN_3043;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_8_state_state <= _GEN_3043;
        end else if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_8_state_state <= _GEN_3043;
        end
      end else begin
        TBEMemory_8_state_state <= _GEN_3043;
      end
    end else begin
      TBEMemory_8_state_state <= _GEN_3557;
    end
    if (reset) begin
      TBEMemory_8_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'h8 == idxAlloc[3:0]) begin
        TBEMemory_8_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h8 == idxAlloc[3:0]) begin
          TBEMemory_8_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEMemory_8_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEMemory_8_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEMemory_8_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEMemory_8_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEMemory_8_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEMemory_8_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEMemory_8_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h8 == idxUpdate_0[3:0]) begin
                        TBEMemory_8_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEMemory_8_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEMemory_8_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h8 == idxUpdate_0[3:0]) begin
                        TBEMemory_8_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h8 == idxAlloc[3:0]) begin
                        TBEMemory_8_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'h8 == idxUpdate_0[3:0]) begin
                        TBEMemory_8_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h8 == idxUpdate_0[3:0]) begin
                          TBEMemory_8_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEMemory_8_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEMemory_8_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h8 == idxUpdate_0[3:0]) begin
                        TBEMemory_8_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_8_way <= _GEN_457;
                end
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEMemory_8_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_8_way <= _GEN_457;
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_way <= 3'h2;
                  end else begin
                    TBEMemory_8_way <= _GEN_457;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_8_way <= _GEN_457;
                  end else if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_8_way <= _GEN_457;
                  end
                end else begin
                  TBEMemory_8_way <= _GEN_457;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEMemory_8_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_8_way <= _GEN_457;
                    end
                  end else if (_T_111) begin
                    if (4'h8 == idxUpdate_1[3:0]) begin
                      TBEMemory_8_way <= 3'h2;
                    end else begin
                      TBEMemory_8_way <= _GEN_457;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_8_way <= _GEN_457;
                    end else if (4'h8 == idxUpdate_1[3:0]) begin
                      TBEMemory_8_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_8_way <= _GEN_457;
                    end
                  end else begin
                    TBEMemory_8_way <= _GEN_457;
                  end
                end else if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEMemory_8_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_8_way <= _GEN_457;
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_way <= 3'h2;
                  end else begin
                    TBEMemory_8_way <= _GEN_457;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_8_way <= _GEN_457;
                  end else if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_8_way <= _GEN_457;
                  end
                end else begin
                  TBEMemory_8_way <= _GEN_457;
                end
              end else begin
                TBEMemory_8_way <= _GEN_971;
              end
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEMemory_8_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_8_way <= _GEN_971;
                end
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_way <= 3'h2;
                end else begin
                  TBEMemory_8_way <= _GEN_971;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_8_way <= _GEN_971;
                end else if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_8_way <= _GEN_971;
                end
              end else begin
                TBEMemory_8_way <= _GEN_971;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEMemory_8_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_8_way <= _GEN_971;
                  end
                end else if (_T_133) begin
                  if (4'h8 == idxUpdate_2[3:0]) begin
                    TBEMemory_8_way <= 3'h2;
                  end else begin
                    TBEMemory_8_way <= _GEN_971;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_8_way <= _GEN_971;
                  end else if (4'h8 == idxUpdate_2[3:0]) begin
                    TBEMemory_8_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_8_way <= _GEN_971;
                  end
                end else begin
                  TBEMemory_8_way <= _GEN_971;
                end
              end else if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEMemory_8_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_8_way <= _GEN_971;
                end
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_way <= 3'h2;
                end else begin
                  TBEMemory_8_way <= _GEN_971;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_8_way <= _GEN_971;
                end else if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_8_way <= _GEN_971;
                end
              end else begin
                TBEMemory_8_way <= _GEN_971;
              end
            end else begin
              TBEMemory_8_way <= _GEN_1485;
            end
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEMemory_8_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_8_way <= _GEN_1485;
              end
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_way <= 3'h2;
              end else begin
                TBEMemory_8_way <= _GEN_1485;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_8_way <= _GEN_1485;
              end else if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_8_way <= _GEN_1485;
              end
            end else begin
              TBEMemory_8_way <= _GEN_1485;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEMemory_8_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_8_way <= _GEN_1485;
                end
              end else if (_T_155) begin
                if (4'h8 == idxUpdate_3[3:0]) begin
                  TBEMemory_8_way <= 3'h2;
                end else begin
                  TBEMemory_8_way <= _GEN_1485;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_8_way <= _GEN_1485;
                end else if (4'h8 == idxUpdate_3[3:0]) begin
                  TBEMemory_8_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_8_way <= _GEN_1485;
                end
              end else begin
                TBEMemory_8_way <= _GEN_1485;
              end
            end else if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEMemory_8_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_8_way <= _GEN_1485;
              end
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_way <= 3'h2;
              end else begin
                TBEMemory_8_way <= _GEN_1485;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_8_way <= _GEN_1485;
              end else if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_8_way <= _GEN_1485;
              end
            end else begin
              TBEMemory_8_way <= _GEN_1485;
            end
          end else begin
            TBEMemory_8_way <= _GEN_1999;
          end
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEMemory_8_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_8_way <= _GEN_1999;
            end
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_way <= 3'h2;
            end else begin
              TBEMemory_8_way <= _GEN_1999;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_8_way <= _GEN_1999;
            end else if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_8_way <= _GEN_1999;
            end
          end else begin
            TBEMemory_8_way <= _GEN_1999;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEMemory_8_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_8_way <= _GEN_1999;
              end
            end else if (_T_177) begin
              if (4'h8 == idxUpdate_4[3:0]) begin
                TBEMemory_8_way <= 3'h2;
              end else begin
                TBEMemory_8_way <= _GEN_1999;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_8_way <= _GEN_1999;
              end else if (4'h8 == idxUpdate_4[3:0]) begin
                TBEMemory_8_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_8_way <= _GEN_1999;
              end
            end else begin
              TBEMemory_8_way <= _GEN_1999;
            end
          end else if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEMemory_8_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_8_way <= _GEN_1999;
            end
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_way <= 3'h2;
            end else begin
              TBEMemory_8_way <= _GEN_1999;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_8_way <= _GEN_1999;
            end else if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_8_way <= _GEN_1999;
            end
          end else begin
            TBEMemory_8_way <= _GEN_1999;
          end
        end else begin
          TBEMemory_8_way <= _GEN_2513;
        end
      end else if (_T_221) begin
        if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEMemory_8_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_8_way <= _GEN_2513;
          end
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_way <= 3'h2;
          end else begin
            TBEMemory_8_way <= _GEN_2513;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_8_way <= _GEN_2513;
          end else if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_8_way <= _GEN_2513;
          end
        end else begin
          TBEMemory_8_way <= _GEN_2513;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEMemory_8_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_8_way <= _GEN_2513;
            end
          end else if (_T_199) begin
            if (4'h8 == idxUpdate_5[3:0]) begin
              TBEMemory_8_way <= 3'h2;
            end else begin
              TBEMemory_8_way <= _GEN_2513;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_8_way <= _GEN_2513;
            end else if (4'h8 == idxUpdate_5[3:0]) begin
              TBEMemory_8_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_8_way <= _GEN_2513;
            end
          end else begin
            TBEMemory_8_way <= _GEN_2513;
          end
        end else if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEMemory_8_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_8_way <= _GEN_2513;
          end
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_way <= 3'h2;
          end else begin
            TBEMemory_8_way <= _GEN_2513;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_8_way <= _GEN_2513;
          end else if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_8_way <= _GEN_2513;
          end
        end else begin
          TBEMemory_8_way <= _GEN_2513;
        end
      end else begin
        TBEMemory_8_way <= _GEN_3027;
      end
    end else if (_T_243) begin
      if (4'h8 == idxUpdate_7[3:0]) begin
        TBEMemory_8_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'h8 == idxAlloc[3:0]) begin
          TBEMemory_8_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_8_way <= _GEN_3027;
        end
      end else if (_T_221) begin
        if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_way <= 3'h2;
        end else begin
          TBEMemory_8_way <= _GEN_3027;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_8_way <= _GEN_3027;
        end else if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_8_way <= _GEN_3027;
        end
      end else begin
        TBEMemory_8_way <= _GEN_3027;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEMemory_8_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_8_way <= _GEN_3027;
          end
        end else if (_T_221) begin
          if (4'h8 == idxUpdate_6[3:0]) begin
            TBEMemory_8_way <= 3'h2;
          end else begin
            TBEMemory_8_way <= _GEN_3027;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_8_way <= _GEN_3027;
          end else if (4'h8 == idxUpdate_6[3:0]) begin
            TBEMemory_8_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_8_way <= _GEN_3027;
          end
        end else begin
          TBEMemory_8_way <= _GEN_3027;
        end
      end else if (4'h8 == idxUpdate_7[3:0]) begin
        TBEMemory_8_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h8 == idxAlloc[3:0]) begin
          TBEMemory_8_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_8_way <= _GEN_3027;
        end
      end else if (_T_221) begin
        if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_way <= 3'h2;
        end else begin
          TBEMemory_8_way <= _GEN_3027;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_8_way <= _GEN_3027;
        end else if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_8_way <= _GEN_3027;
        end
      end else begin
        TBEMemory_8_way <= _GEN_3027;
      end
    end else begin
      TBEMemory_8_way <= _GEN_3541;
    end
    if (reset) begin
      TBEMemory_8_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h8 == idxAlloc[3:0]) begin
        TBEMemory_8_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'h8 == idxAlloc[3:0]) begin
          TBEMemory_8_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEMemory_8_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEMemory_8_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEMemory_8_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEMemory_8_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEMemory_8_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEMemory_8_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEMemory_8_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h8 == idxUpdate_0[3:0]) begin
                        TBEMemory_8_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEMemory_8_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEMemory_8_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h8 == idxUpdate_0[3:0]) begin
                        TBEMemory_8_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h8 == idxUpdate_1[3:0]) begin
                      TBEMemory_8_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'h8 == idxAlloc[3:0]) begin
                        TBEMemory_8_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'h8 == idxUpdate_0[3:0]) begin
                        TBEMemory_8_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'h8 == idxUpdate_0[3:0]) begin
                          TBEMemory_8_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEMemory_8_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEMemory_8_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h8 == idxUpdate_0[3:0]) begin
                        TBEMemory_8_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_441;
                end
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEMemory_8_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_441;
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_441;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h8 == idxUpdate_1[3:0]) begin
                      TBEMemory_8_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_8_fields_0 <= _GEN_441;
                    end
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_441;
                  end
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_441;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h8 == idxUpdate_2[3:0]) begin
                    TBEMemory_8_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEMemory_8_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_8_fields_0 <= _GEN_441;
                    end
                  end else if (_T_111) begin
                    if (4'h8 == idxUpdate_1[3:0]) begin
                      TBEMemory_8_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_8_fields_0 <= _GEN_441;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'h8 == idxUpdate_1[3:0]) begin
                        TBEMemory_8_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_8_fields_0 <= _GEN_441;
                      end
                    end else begin
                      TBEMemory_8_fields_0 <= _GEN_441;
                    end
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_441;
                  end
                end else if (isAlloc_1) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEMemory_8_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_441;
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEMemory_8_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_441;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h8 == idxUpdate_1[3:0]) begin
                      TBEMemory_8_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_8_fields_0 <= _GEN_441;
                    end
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_441;
                  end
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_441;
                end
              end else begin
                TBEMemory_8_fields_0 <= _GEN_955;
              end
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEMemory_8_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_955;
                end
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_955;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h8 == idxUpdate_2[3:0]) begin
                    TBEMemory_8_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_955;
                  end
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_955;
                end
              end else begin
                TBEMemory_8_fields_0 <= _GEN_955;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h8 == idxUpdate_3[3:0]) begin
                  TBEMemory_8_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEMemory_8_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_955;
                  end
                end else if (_T_133) begin
                  if (4'h8 == idxUpdate_2[3:0]) begin
                    TBEMemory_8_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_955;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'h8 == idxUpdate_2[3:0]) begin
                      TBEMemory_8_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_8_fields_0 <= _GEN_955;
                    end
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_955;
                  end
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_955;
                end
              end else if (isAlloc_2) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEMemory_8_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_955;
                end
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEMemory_8_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_955;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h8 == idxUpdate_2[3:0]) begin
                    TBEMemory_8_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_955;
                  end
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_955;
                end
              end else begin
                TBEMemory_8_fields_0 <= _GEN_955;
              end
            end else begin
              TBEMemory_8_fields_0 <= _GEN_1469;
            end
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEMemory_8_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_8_fields_0 <= _GEN_1469;
              end
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_fields_0 <= 32'h0;
              end else begin
                TBEMemory_8_fields_0 <= _GEN_1469;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h8 == idxUpdate_3[3:0]) begin
                  TBEMemory_8_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_1469;
                end
              end else begin
                TBEMemory_8_fields_0 <= _GEN_1469;
              end
            end else begin
              TBEMemory_8_fields_0 <= _GEN_1469;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h8 == idxUpdate_4[3:0]) begin
                TBEMemory_8_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEMemory_8_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_1469;
                end
              end else if (_T_155) begin
                if (4'h8 == idxUpdate_3[3:0]) begin
                  TBEMemory_8_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_1469;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'h8 == idxUpdate_3[3:0]) begin
                    TBEMemory_8_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_8_fields_0 <= _GEN_1469;
                  end
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_1469;
                end
              end else begin
                TBEMemory_8_fields_0 <= _GEN_1469;
              end
            end else if (isAlloc_3) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEMemory_8_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_8_fields_0 <= _GEN_1469;
              end
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEMemory_8_fields_0 <= 32'h0;
              end else begin
                TBEMemory_8_fields_0 <= _GEN_1469;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h8 == idxUpdate_3[3:0]) begin
                  TBEMemory_8_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_1469;
                end
              end else begin
                TBEMemory_8_fields_0 <= _GEN_1469;
              end
            end else begin
              TBEMemory_8_fields_0 <= _GEN_1469;
            end
          end else begin
            TBEMemory_8_fields_0 <= _GEN_1983;
          end
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEMemory_8_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_8_fields_0 <= _GEN_1983;
            end
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_fields_0 <= 32'h0;
            end else begin
              TBEMemory_8_fields_0 <= _GEN_1983;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h8 == idxUpdate_4[3:0]) begin
                TBEMemory_8_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_8_fields_0 <= _GEN_1983;
              end
            end else begin
              TBEMemory_8_fields_0 <= _GEN_1983;
            end
          end else begin
            TBEMemory_8_fields_0 <= _GEN_1983;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h8 == idxUpdate_5[3:0]) begin
              TBEMemory_8_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEMemory_8_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_8_fields_0 <= _GEN_1983;
              end
            end else if (_T_177) begin
              if (4'h8 == idxUpdate_4[3:0]) begin
                TBEMemory_8_fields_0 <= 32'h0;
              end else begin
                TBEMemory_8_fields_0 <= _GEN_1983;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'h8 == idxUpdate_4[3:0]) begin
                  TBEMemory_8_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_8_fields_0 <= _GEN_1983;
                end
              end else begin
                TBEMemory_8_fields_0 <= _GEN_1983;
              end
            end else begin
              TBEMemory_8_fields_0 <= _GEN_1983;
            end
          end else if (isAlloc_4) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEMemory_8_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_8_fields_0 <= _GEN_1983;
            end
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEMemory_8_fields_0 <= 32'h0;
            end else begin
              TBEMemory_8_fields_0 <= _GEN_1983;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h8 == idxUpdate_4[3:0]) begin
                TBEMemory_8_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_8_fields_0 <= _GEN_1983;
              end
            end else begin
              TBEMemory_8_fields_0 <= _GEN_1983;
            end
          end else begin
            TBEMemory_8_fields_0 <= _GEN_1983;
          end
        end else begin
          TBEMemory_8_fields_0 <= _GEN_2497;
        end
      end else if (_T_221) begin
        if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEMemory_8_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_8_fields_0 <= _GEN_2497;
          end
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_fields_0 <= 32'h0;
          end else begin
            TBEMemory_8_fields_0 <= _GEN_2497;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h8 == idxUpdate_5[3:0]) begin
              TBEMemory_8_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_8_fields_0 <= _GEN_2497;
            end
          end else begin
            TBEMemory_8_fields_0 <= _GEN_2497;
          end
        end else begin
          TBEMemory_8_fields_0 <= _GEN_2497;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h8 == idxUpdate_6[3:0]) begin
            TBEMemory_8_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEMemory_8_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_8_fields_0 <= _GEN_2497;
            end
          end else if (_T_199) begin
            if (4'h8 == idxUpdate_5[3:0]) begin
              TBEMemory_8_fields_0 <= 32'h0;
            end else begin
              TBEMemory_8_fields_0 <= _GEN_2497;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'h8 == idxUpdate_5[3:0]) begin
                TBEMemory_8_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_8_fields_0 <= _GEN_2497;
              end
            end else begin
              TBEMemory_8_fields_0 <= _GEN_2497;
            end
          end else begin
            TBEMemory_8_fields_0 <= _GEN_2497;
          end
        end else if (isAlloc_5) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEMemory_8_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_8_fields_0 <= _GEN_2497;
          end
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEMemory_8_fields_0 <= 32'h0;
          end else begin
            TBEMemory_8_fields_0 <= _GEN_2497;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h8 == idxUpdate_5[3:0]) begin
              TBEMemory_8_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_8_fields_0 <= _GEN_2497;
            end
          end else begin
            TBEMemory_8_fields_0 <= _GEN_2497;
          end
        end else begin
          TBEMemory_8_fields_0 <= _GEN_2497;
        end
      end else begin
        TBEMemory_8_fields_0 <= _GEN_3011;
      end
    end else if (_T_243) begin
      if (4'h8 == idxUpdate_7[3:0]) begin
        TBEMemory_8_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h8 == idxAlloc[3:0]) begin
          TBEMemory_8_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_8_fields_0 <= _GEN_3011;
        end
      end else if (_T_221) begin
        if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_fields_0 <= 32'h0;
        end else begin
          TBEMemory_8_fields_0 <= _GEN_3011;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h8 == idxUpdate_6[3:0]) begin
            TBEMemory_8_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_8_fields_0 <= _GEN_3011;
          end
        end else begin
          TBEMemory_8_fields_0 <= _GEN_3011;
        end
      end else begin
        TBEMemory_8_fields_0 <= _GEN_3011;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'h8 == idxUpdate_7[3:0]) begin
          TBEMemory_8_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEMemory_8_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_8_fields_0 <= _GEN_3011;
          end
        end else if (_T_221) begin
          if (4'h8 == idxUpdate_6[3:0]) begin
            TBEMemory_8_fields_0 <= 32'h0;
          end else begin
            TBEMemory_8_fields_0 <= _GEN_3011;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'h8 == idxUpdate_6[3:0]) begin
              TBEMemory_8_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_8_fields_0 <= _GEN_3011;
            end
          end else begin
            TBEMemory_8_fields_0 <= _GEN_3011;
          end
        end else begin
          TBEMemory_8_fields_0 <= _GEN_3011;
        end
      end else if (isAlloc_6) begin
        if (4'h8 == idxAlloc[3:0]) begin
          TBEMemory_8_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_8_fields_0 <= _GEN_3011;
        end
      end else if (_T_221) begin
        if (4'h8 == idxUpdate_6[3:0]) begin
          TBEMemory_8_fields_0 <= 32'h0;
        end else begin
          TBEMemory_8_fields_0 <= _GEN_3011;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h8 == idxUpdate_6[3:0]) begin
            TBEMemory_8_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_8_fields_0 <= _GEN_3011;
          end
        end else begin
          TBEMemory_8_fields_0 <= _GEN_3011;
        end
      end else begin
        TBEMemory_8_fields_0 <= _GEN_3011;
      end
    end else begin
      TBEMemory_8_fields_0 <= _GEN_3525;
    end
    if (reset) begin
      TBEMemory_9_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'h9 == idxAlloc[3:0]) begin
        TBEMemory_9_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h9 == idxAlloc[3:0]) begin
          TBEMemory_9_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEMemory_9_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEMemory_9_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEMemory_9_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEMemory_9_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEMemory_9_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEMemory_9_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEMemory_9_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h9 == idxUpdate_0[3:0]) begin
                        TBEMemory_9_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEMemory_9_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEMemory_9_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h9 == idxUpdate_0[3:0]) begin
                        TBEMemory_9_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h9 == idxAlloc[3:0]) begin
                        TBEMemory_9_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'h9 == idxUpdate_0[3:0]) begin
                        TBEMemory_9_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h9 == idxUpdate_0[3:0]) begin
                          TBEMemory_9_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEMemory_9_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEMemory_9_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h9 == idxUpdate_0[3:0]) begin
                        TBEMemory_9_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_9_state_state <= _GEN_474;
                end
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEMemory_9_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_9_state_state <= _GEN_474;
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_state_state <= 2'h0;
                  end else begin
                    TBEMemory_9_state_state <= _GEN_474;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_9_state_state <= _GEN_474;
                  end else if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_9_state_state <= _GEN_474;
                  end
                end else begin
                  TBEMemory_9_state_state <= _GEN_474;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEMemory_9_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_9_state_state <= _GEN_474;
                    end
                  end else if (_T_111) begin
                    if (4'h9 == idxUpdate_1[3:0]) begin
                      TBEMemory_9_state_state <= 2'h0;
                    end else begin
                      TBEMemory_9_state_state <= _GEN_474;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_9_state_state <= _GEN_474;
                    end else if (4'h9 == idxUpdate_1[3:0]) begin
                      TBEMemory_9_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_9_state_state <= _GEN_474;
                    end
                  end else begin
                    TBEMemory_9_state_state <= _GEN_474;
                  end
                end else if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEMemory_9_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_9_state_state <= _GEN_474;
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_state_state <= 2'h0;
                  end else begin
                    TBEMemory_9_state_state <= _GEN_474;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_9_state_state <= _GEN_474;
                  end else if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_9_state_state <= _GEN_474;
                  end
                end else begin
                  TBEMemory_9_state_state <= _GEN_474;
                end
              end else begin
                TBEMemory_9_state_state <= _GEN_988;
              end
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEMemory_9_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_9_state_state <= _GEN_988;
                end
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_state_state <= 2'h0;
                end else begin
                  TBEMemory_9_state_state <= _GEN_988;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_9_state_state <= _GEN_988;
                end else if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_9_state_state <= _GEN_988;
                end
              end else begin
                TBEMemory_9_state_state <= _GEN_988;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEMemory_9_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_9_state_state <= _GEN_988;
                  end
                end else if (_T_133) begin
                  if (4'h9 == idxUpdate_2[3:0]) begin
                    TBEMemory_9_state_state <= 2'h0;
                  end else begin
                    TBEMemory_9_state_state <= _GEN_988;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_9_state_state <= _GEN_988;
                  end else if (4'h9 == idxUpdate_2[3:0]) begin
                    TBEMemory_9_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_9_state_state <= _GEN_988;
                  end
                end else begin
                  TBEMemory_9_state_state <= _GEN_988;
                end
              end else if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEMemory_9_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_9_state_state <= _GEN_988;
                end
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_state_state <= 2'h0;
                end else begin
                  TBEMemory_9_state_state <= _GEN_988;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_9_state_state <= _GEN_988;
                end else if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_9_state_state <= _GEN_988;
                end
              end else begin
                TBEMemory_9_state_state <= _GEN_988;
              end
            end else begin
              TBEMemory_9_state_state <= _GEN_1502;
            end
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEMemory_9_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_9_state_state <= _GEN_1502;
              end
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_state_state <= 2'h0;
              end else begin
                TBEMemory_9_state_state <= _GEN_1502;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_9_state_state <= _GEN_1502;
              end else if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_9_state_state <= _GEN_1502;
              end
            end else begin
              TBEMemory_9_state_state <= _GEN_1502;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEMemory_9_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_9_state_state <= _GEN_1502;
                end
              end else if (_T_155) begin
                if (4'h9 == idxUpdate_3[3:0]) begin
                  TBEMemory_9_state_state <= 2'h0;
                end else begin
                  TBEMemory_9_state_state <= _GEN_1502;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_9_state_state <= _GEN_1502;
                end else if (4'h9 == idxUpdate_3[3:0]) begin
                  TBEMemory_9_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_9_state_state <= _GEN_1502;
                end
              end else begin
                TBEMemory_9_state_state <= _GEN_1502;
              end
            end else if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEMemory_9_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_9_state_state <= _GEN_1502;
              end
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_state_state <= 2'h0;
              end else begin
                TBEMemory_9_state_state <= _GEN_1502;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_9_state_state <= _GEN_1502;
              end else if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_9_state_state <= _GEN_1502;
              end
            end else begin
              TBEMemory_9_state_state <= _GEN_1502;
            end
          end else begin
            TBEMemory_9_state_state <= _GEN_2016;
          end
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEMemory_9_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_9_state_state <= _GEN_2016;
            end
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_state_state <= 2'h0;
            end else begin
              TBEMemory_9_state_state <= _GEN_2016;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_9_state_state <= _GEN_2016;
            end else if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_9_state_state <= _GEN_2016;
            end
          end else begin
            TBEMemory_9_state_state <= _GEN_2016;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEMemory_9_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_9_state_state <= _GEN_2016;
              end
            end else if (_T_177) begin
              if (4'h9 == idxUpdate_4[3:0]) begin
                TBEMemory_9_state_state <= 2'h0;
              end else begin
                TBEMemory_9_state_state <= _GEN_2016;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_9_state_state <= _GEN_2016;
              end else if (4'h9 == idxUpdate_4[3:0]) begin
                TBEMemory_9_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_9_state_state <= _GEN_2016;
              end
            end else begin
              TBEMemory_9_state_state <= _GEN_2016;
            end
          end else if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEMemory_9_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_9_state_state <= _GEN_2016;
            end
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_state_state <= 2'h0;
            end else begin
              TBEMemory_9_state_state <= _GEN_2016;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_9_state_state <= _GEN_2016;
            end else if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_9_state_state <= _GEN_2016;
            end
          end else begin
            TBEMemory_9_state_state <= _GEN_2016;
          end
        end else begin
          TBEMemory_9_state_state <= _GEN_2530;
        end
      end else if (_T_221) begin
        if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEMemory_9_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_9_state_state <= _GEN_2530;
          end
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_state_state <= 2'h0;
          end else begin
            TBEMemory_9_state_state <= _GEN_2530;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_9_state_state <= _GEN_2530;
          end else if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_9_state_state <= _GEN_2530;
          end
        end else begin
          TBEMemory_9_state_state <= _GEN_2530;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEMemory_9_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_9_state_state <= _GEN_2530;
            end
          end else if (_T_199) begin
            if (4'h9 == idxUpdate_5[3:0]) begin
              TBEMemory_9_state_state <= 2'h0;
            end else begin
              TBEMemory_9_state_state <= _GEN_2530;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_9_state_state <= _GEN_2530;
            end else if (4'h9 == idxUpdate_5[3:0]) begin
              TBEMemory_9_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_9_state_state <= _GEN_2530;
            end
          end else begin
            TBEMemory_9_state_state <= _GEN_2530;
          end
        end else if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEMemory_9_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_9_state_state <= _GEN_2530;
          end
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_state_state <= 2'h0;
          end else begin
            TBEMemory_9_state_state <= _GEN_2530;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_9_state_state <= _GEN_2530;
          end else if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_9_state_state <= _GEN_2530;
          end
        end else begin
          TBEMemory_9_state_state <= _GEN_2530;
        end
      end else begin
        TBEMemory_9_state_state <= _GEN_3044;
      end
    end else if (_T_243) begin
      if (4'h9 == idxUpdate_7[3:0]) begin
        TBEMemory_9_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'h9 == idxAlloc[3:0]) begin
          TBEMemory_9_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_9_state_state <= _GEN_3044;
        end
      end else if (_T_221) begin
        if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_state_state <= 2'h0;
        end else begin
          TBEMemory_9_state_state <= _GEN_3044;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_9_state_state <= _GEN_3044;
        end else if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_9_state_state <= _GEN_3044;
        end
      end else begin
        TBEMemory_9_state_state <= _GEN_3044;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEMemory_9_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_9_state_state <= _GEN_3044;
          end
        end else if (_T_221) begin
          if (4'h9 == idxUpdate_6[3:0]) begin
            TBEMemory_9_state_state <= 2'h0;
          end else begin
            TBEMemory_9_state_state <= _GEN_3044;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_9_state_state <= _GEN_3044;
          end else if (4'h9 == idxUpdate_6[3:0]) begin
            TBEMemory_9_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_9_state_state <= _GEN_3044;
          end
        end else begin
          TBEMemory_9_state_state <= _GEN_3044;
        end
      end else if (4'h9 == idxUpdate_7[3:0]) begin
        TBEMemory_9_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'h9 == idxAlloc[3:0]) begin
          TBEMemory_9_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_9_state_state <= _GEN_3044;
        end
      end else if (_T_221) begin
        if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_state_state <= 2'h0;
        end else begin
          TBEMemory_9_state_state <= _GEN_3044;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_9_state_state <= _GEN_3044;
        end else if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_9_state_state <= _GEN_3044;
        end
      end else begin
        TBEMemory_9_state_state <= _GEN_3044;
      end
    end else begin
      TBEMemory_9_state_state <= _GEN_3558;
    end
    if (reset) begin
      TBEMemory_9_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'h9 == idxAlloc[3:0]) begin
        TBEMemory_9_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h9 == idxAlloc[3:0]) begin
          TBEMemory_9_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEMemory_9_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEMemory_9_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEMemory_9_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEMemory_9_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEMemory_9_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEMemory_9_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEMemory_9_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h9 == idxUpdate_0[3:0]) begin
                        TBEMemory_9_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEMemory_9_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEMemory_9_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h9 == idxUpdate_0[3:0]) begin
                        TBEMemory_9_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'h9 == idxAlloc[3:0]) begin
                        TBEMemory_9_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'h9 == idxUpdate_0[3:0]) begin
                        TBEMemory_9_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'h9 == idxUpdate_0[3:0]) begin
                          TBEMemory_9_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEMemory_9_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEMemory_9_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'h9 == idxUpdate_0[3:0]) begin
                        TBEMemory_9_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_9_way <= _GEN_458;
                end
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEMemory_9_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_9_way <= _GEN_458;
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_way <= 3'h2;
                  end else begin
                    TBEMemory_9_way <= _GEN_458;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_9_way <= _GEN_458;
                  end else if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_9_way <= _GEN_458;
                  end
                end else begin
                  TBEMemory_9_way <= _GEN_458;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEMemory_9_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_9_way <= _GEN_458;
                    end
                  end else if (_T_111) begin
                    if (4'h9 == idxUpdate_1[3:0]) begin
                      TBEMemory_9_way <= 3'h2;
                    end else begin
                      TBEMemory_9_way <= _GEN_458;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_9_way <= _GEN_458;
                    end else if (4'h9 == idxUpdate_1[3:0]) begin
                      TBEMemory_9_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_9_way <= _GEN_458;
                    end
                  end else begin
                    TBEMemory_9_way <= _GEN_458;
                  end
                end else if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEMemory_9_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_9_way <= _GEN_458;
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_way <= 3'h2;
                  end else begin
                    TBEMemory_9_way <= _GEN_458;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_9_way <= _GEN_458;
                  end else if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_9_way <= _GEN_458;
                  end
                end else begin
                  TBEMemory_9_way <= _GEN_458;
                end
              end else begin
                TBEMemory_9_way <= _GEN_972;
              end
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEMemory_9_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_9_way <= _GEN_972;
                end
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_way <= 3'h2;
                end else begin
                  TBEMemory_9_way <= _GEN_972;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_9_way <= _GEN_972;
                end else if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_9_way <= _GEN_972;
                end
              end else begin
                TBEMemory_9_way <= _GEN_972;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEMemory_9_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_9_way <= _GEN_972;
                  end
                end else if (_T_133) begin
                  if (4'h9 == idxUpdate_2[3:0]) begin
                    TBEMemory_9_way <= 3'h2;
                  end else begin
                    TBEMemory_9_way <= _GEN_972;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_9_way <= _GEN_972;
                  end else if (4'h9 == idxUpdate_2[3:0]) begin
                    TBEMemory_9_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_9_way <= _GEN_972;
                  end
                end else begin
                  TBEMemory_9_way <= _GEN_972;
                end
              end else if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEMemory_9_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_9_way <= _GEN_972;
                end
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_way <= 3'h2;
                end else begin
                  TBEMemory_9_way <= _GEN_972;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_9_way <= _GEN_972;
                end else if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_9_way <= _GEN_972;
                end
              end else begin
                TBEMemory_9_way <= _GEN_972;
              end
            end else begin
              TBEMemory_9_way <= _GEN_1486;
            end
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEMemory_9_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_9_way <= _GEN_1486;
              end
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_way <= 3'h2;
              end else begin
                TBEMemory_9_way <= _GEN_1486;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_9_way <= _GEN_1486;
              end else if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_9_way <= _GEN_1486;
              end
            end else begin
              TBEMemory_9_way <= _GEN_1486;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEMemory_9_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_9_way <= _GEN_1486;
                end
              end else if (_T_155) begin
                if (4'h9 == idxUpdate_3[3:0]) begin
                  TBEMemory_9_way <= 3'h2;
                end else begin
                  TBEMemory_9_way <= _GEN_1486;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_9_way <= _GEN_1486;
                end else if (4'h9 == idxUpdate_3[3:0]) begin
                  TBEMemory_9_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_9_way <= _GEN_1486;
                end
              end else begin
                TBEMemory_9_way <= _GEN_1486;
              end
            end else if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEMemory_9_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_9_way <= _GEN_1486;
              end
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_way <= 3'h2;
              end else begin
                TBEMemory_9_way <= _GEN_1486;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_9_way <= _GEN_1486;
              end else if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_9_way <= _GEN_1486;
              end
            end else begin
              TBEMemory_9_way <= _GEN_1486;
            end
          end else begin
            TBEMemory_9_way <= _GEN_2000;
          end
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEMemory_9_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_9_way <= _GEN_2000;
            end
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_way <= 3'h2;
            end else begin
              TBEMemory_9_way <= _GEN_2000;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_9_way <= _GEN_2000;
            end else if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_9_way <= _GEN_2000;
            end
          end else begin
            TBEMemory_9_way <= _GEN_2000;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEMemory_9_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_9_way <= _GEN_2000;
              end
            end else if (_T_177) begin
              if (4'h9 == idxUpdate_4[3:0]) begin
                TBEMemory_9_way <= 3'h2;
              end else begin
                TBEMemory_9_way <= _GEN_2000;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_9_way <= _GEN_2000;
              end else if (4'h9 == idxUpdate_4[3:0]) begin
                TBEMemory_9_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_9_way <= _GEN_2000;
              end
            end else begin
              TBEMemory_9_way <= _GEN_2000;
            end
          end else if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEMemory_9_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_9_way <= _GEN_2000;
            end
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_way <= 3'h2;
            end else begin
              TBEMemory_9_way <= _GEN_2000;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_9_way <= _GEN_2000;
            end else if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_9_way <= _GEN_2000;
            end
          end else begin
            TBEMemory_9_way <= _GEN_2000;
          end
        end else begin
          TBEMemory_9_way <= _GEN_2514;
        end
      end else if (_T_221) begin
        if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEMemory_9_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_9_way <= _GEN_2514;
          end
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_way <= 3'h2;
          end else begin
            TBEMemory_9_way <= _GEN_2514;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_9_way <= _GEN_2514;
          end else if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_9_way <= _GEN_2514;
          end
        end else begin
          TBEMemory_9_way <= _GEN_2514;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEMemory_9_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_9_way <= _GEN_2514;
            end
          end else if (_T_199) begin
            if (4'h9 == idxUpdate_5[3:0]) begin
              TBEMemory_9_way <= 3'h2;
            end else begin
              TBEMemory_9_way <= _GEN_2514;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_9_way <= _GEN_2514;
            end else if (4'h9 == idxUpdate_5[3:0]) begin
              TBEMemory_9_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_9_way <= _GEN_2514;
            end
          end else begin
            TBEMemory_9_way <= _GEN_2514;
          end
        end else if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEMemory_9_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_9_way <= _GEN_2514;
          end
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_way <= 3'h2;
          end else begin
            TBEMemory_9_way <= _GEN_2514;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_9_way <= _GEN_2514;
          end else if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_9_way <= _GEN_2514;
          end
        end else begin
          TBEMemory_9_way <= _GEN_2514;
        end
      end else begin
        TBEMemory_9_way <= _GEN_3028;
      end
    end else if (_T_243) begin
      if (4'h9 == idxUpdate_7[3:0]) begin
        TBEMemory_9_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'h9 == idxAlloc[3:0]) begin
          TBEMemory_9_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_9_way <= _GEN_3028;
        end
      end else if (_T_221) begin
        if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_way <= 3'h2;
        end else begin
          TBEMemory_9_way <= _GEN_3028;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_9_way <= _GEN_3028;
        end else if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_9_way <= _GEN_3028;
        end
      end else begin
        TBEMemory_9_way <= _GEN_3028;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEMemory_9_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_9_way <= _GEN_3028;
          end
        end else if (_T_221) begin
          if (4'h9 == idxUpdate_6[3:0]) begin
            TBEMemory_9_way <= 3'h2;
          end else begin
            TBEMemory_9_way <= _GEN_3028;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_9_way <= _GEN_3028;
          end else if (4'h9 == idxUpdate_6[3:0]) begin
            TBEMemory_9_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_9_way <= _GEN_3028;
          end
        end else begin
          TBEMemory_9_way <= _GEN_3028;
        end
      end else if (4'h9 == idxUpdate_7[3:0]) begin
        TBEMemory_9_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'h9 == idxAlloc[3:0]) begin
          TBEMemory_9_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_9_way <= _GEN_3028;
        end
      end else if (_T_221) begin
        if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_way <= 3'h2;
        end else begin
          TBEMemory_9_way <= _GEN_3028;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_9_way <= _GEN_3028;
        end else if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_9_way <= _GEN_3028;
        end
      end else begin
        TBEMemory_9_way <= _GEN_3028;
      end
    end else begin
      TBEMemory_9_way <= _GEN_3542;
    end
    if (reset) begin
      TBEMemory_9_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h9 == idxAlloc[3:0]) begin
        TBEMemory_9_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'h9 == idxAlloc[3:0]) begin
          TBEMemory_9_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEMemory_9_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEMemory_9_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEMemory_9_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEMemory_9_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEMemory_9_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEMemory_9_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEMemory_9_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h9 == idxUpdate_0[3:0]) begin
                        TBEMemory_9_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEMemory_9_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEMemory_9_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h9 == idxUpdate_0[3:0]) begin
                        TBEMemory_9_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h9 == idxUpdate_1[3:0]) begin
                      TBEMemory_9_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'h9 == idxAlloc[3:0]) begin
                        TBEMemory_9_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'h9 == idxUpdate_0[3:0]) begin
                        TBEMemory_9_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'h9 == idxUpdate_0[3:0]) begin
                          TBEMemory_9_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEMemory_9_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEMemory_9_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'h9 == idxUpdate_0[3:0]) begin
                        TBEMemory_9_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_442;
                end
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEMemory_9_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_442;
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_442;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h9 == idxUpdate_1[3:0]) begin
                      TBEMemory_9_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_9_fields_0 <= _GEN_442;
                    end
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_442;
                  end
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_442;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h9 == idxUpdate_2[3:0]) begin
                    TBEMemory_9_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEMemory_9_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_9_fields_0 <= _GEN_442;
                    end
                  end else if (_T_111) begin
                    if (4'h9 == idxUpdate_1[3:0]) begin
                      TBEMemory_9_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_9_fields_0 <= _GEN_442;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'h9 == idxUpdate_1[3:0]) begin
                        TBEMemory_9_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_9_fields_0 <= _GEN_442;
                      end
                    end else begin
                      TBEMemory_9_fields_0 <= _GEN_442;
                    end
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_442;
                  end
                end else if (isAlloc_1) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEMemory_9_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_442;
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEMemory_9_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_442;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'h9 == idxUpdate_1[3:0]) begin
                      TBEMemory_9_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_9_fields_0 <= _GEN_442;
                    end
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_442;
                  end
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_442;
                end
              end else begin
                TBEMemory_9_fields_0 <= _GEN_956;
              end
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEMemory_9_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_956;
                end
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_956;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h9 == idxUpdate_2[3:0]) begin
                    TBEMemory_9_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_956;
                  end
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_956;
                end
              end else begin
                TBEMemory_9_fields_0 <= _GEN_956;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h9 == idxUpdate_3[3:0]) begin
                  TBEMemory_9_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEMemory_9_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_956;
                  end
                end else if (_T_133) begin
                  if (4'h9 == idxUpdate_2[3:0]) begin
                    TBEMemory_9_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_956;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'h9 == idxUpdate_2[3:0]) begin
                      TBEMemory_9_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_9_fields_0 <= _GEN_956;
                    end
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_956;
                  end
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_956;
                end
              end else if (isAlloc_2) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEMemory_9_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_956;
                end
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEMemory_9_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_956;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'h9 == idxUpdate_2[3:0]) begin
                    TBEMemory_9_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_956;
                  end
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_956;
                end
              end else begin
                TBEMemory_9_fields_0 <= _GEN_956;
              end
            end else begin
              TBEMemory_9_fields_0 <= _GEN_1470;
            end
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEMemory_9_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_9_fields_0 <= _GEN_1470;
              end
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_fields_0 <= 32'h0;
              end else begin
                TBEMemory_9_fields_0 <= _GEN_1470;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h9 == idxUpdate_3[3:0]) begin
                  TBEMemory_9_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_1470;
                end
              end else begin
                TBEMemory_9_fields_0 <= _GEN_1470;
              end
            end else begin
              TBEMemory_9_fields_0 <= _GEN_1470;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h9 == idxUpdate_4[3:0]) begin
                TBEMemory_9_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEMemory_9_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_1470;
                end
              end else if (_T_155) begin
                if (4'h9 == idxUpdate_3[3:0]) begin
                  TBEMemory_9_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_1470;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'h9 == idxUpdate_3[3:0]) begin
                    TBEMemory_9_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_9_fields_0 <= _GEN_1470;
                  end
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_1470;
                end
              end else begin
                TBEMemory_9_fields_0 <= _GEN_1470;
              end
            end else if (isAlloc_3) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEMemory_9_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_9_fields_0 <= _GEN_1470;
              end
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEMemory_9_fields_0 <= 32'h0;
              end else begin
                TBEMemory_9_fields_0 <= _GEN_1470;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'h9 == idxUpdate_3[3:0]) begin
                  TBEMemory_9_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_1470;
                end
              end else begin
                TBEMemory_9_fields_0 <= _GEN_1470;
              end
            end else begin
              TBEMemory_9_fields_0 <= _GEN_1470;
            end
          end else begin
            TBEMemory_9_fields_0 <= _GEN_1984;
          end
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEMemory_9_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_9_fields_0 <= _GEN_1984;
            end
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_fields_0 <= 32'h0;
            end else begin
              TBEMemory_9_fields_0 <= _GEN_1984;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h9 == idxUpdate_4[3:0]) begin
                TBEMemory_9_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_9_fields_0 <= _GEN_1984;
              end
            end else begin
              TBEMemory_9_fields_0 <= _GEN_1984;
            end
          end else begin
            TBEMemory_9_fields_0 <= _GEN_1984;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h9 == idxUpdate_5[3:0]) begin
              TBEMemory_9_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEMemory_9_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_9_fields_0 <= _GEN_1984;
              end
            end else if (_T_177) begin
              if (4'h9 == idxUpdate_4[3:0]) begin
                TBEMemory_9_fields_0 <= 32'h0;
              end else begin
                TBEMemory_9_fields_0 <= _GEN_1984;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'h9 == idxUpdate_4[3:0]) begin
                  TBEMemory_9_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_9_fields_0 <= _GEN_1984;
                end
              end else begin
                TBEMemory_9_fields_0 <= _GEN_1984;
              end
            end else begin
              TBEMemory_9_fields_0 <= _GEN_1984;
            end
          end else if (isAlloc_4) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEMemory_9_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_9_fields_0 <= _GEN_1984;
            end
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEMemory_9_fields_0 <= 32'h0;
            end else begin
              TBEMemory_9_fields_0 <= _GEN_1984;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'h9 == idxUpdate_4[3:0]) begin
                TBEMemory_9_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_9_fields_0 <= _GEN_1984;
              end
            end else begin
              TBEMemory_9_fields_0 <= _GEN_1984;
            end
          end else begin
            TBEMemory_9_fields_0 <= _GEN_1984;
          end
        end else begin
          TBEMemory_9_fields_0 <= _GEN_2498;
        end
      end else if (_T_221) begin
        if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEMemory_9_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_9_fields_0 <= _GEN_2498;
          end
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_fields_0 <= 32'h0;
          end else begin
            TBEMemory_9_fields_0 <= _GEN_2498;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h9 == idxUpdate_5[3:0]) begin
              TBEMemory_9_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_9_fields_0 <= _GEN_2498;
            end
          end else begin
            TBEMemory_9_fields_0 <= _GEN_2498;
          end
        end else begin
          TBEMemory_9_fields_0 <= _GEN_2498;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h9 == idxUpdate_6[3:0]) begin
            TBEMemory_9_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEMemory_9_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_9_fields_0 <= _GEN_2498;
            end
          end else if (_T_199) begin
            if (4'h9 == idxUpdate_5[3:0]) begin
              TBEMemory_9_fields_0 <= 32'h0;
            end else begin
              TBEMemory_9_fields_0 <= _GEN_2498;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'h9 == idxUpdate_5[3:0]) begin
                TBEMemory_9_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_9_fields_0 <= _GEN_2498;
              end
            end else begin
              TBEMemory_9_fields_0 <= _GEN_2498;
            end
          end else begin
            TBEMemory_9_fields_0 <= _GEN_2498;
          end
        end else if (isAlloc_5) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEMemory_9_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_9_fields_0 <= _GEN_2498;
          end
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEMemory_9_fields_0 <= 32'h0;
          end else begin
            TBEMemory_9_fields_0 <= _GEN_2498;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'h9 == idxUpdate_5[3:0]) begin
              TBEMemory_9_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_9_fields_0 <= _GEN_2498;
            end
          end else begin
            TBEMemory_9_fields_0 <= _GEN_2498;
          end
        end else begin
          TBEMemory_9_fields_0 <= _GEN_2498;
        end
      end else begin
        TBEMemory_9_fields_0 <= _GEN_3012;
      end
    end else if (_T_243) begin
      if (4'h9 == idxUpdate_7[3:0]) begin
        TBEMemory_9_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h9 == idxAlloc[3:0]) begin
          TBEMemory_9_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_9_fields_0 <= _GEN_3012;
        end
      end else if (_T_221) begin
        if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_fields_0 <= 32'h0;
        end else begin
          TBEMemory_9_fields_0 <= _GEN_3012;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h9 == idxUpdate_6[3:0]) begin
            TBEMemory_9_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_9_fields_0 <= _GEN_3012;
          end
        end else begin
          TBEMemory_9_fields_0 <= _GEN_3012;
        end
      end else begin
        TBEMemory_9_fields_0 <= _GEN_3012;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'h9 == idxUpdate_7[3:0]) begin
          TBEMemory_9_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEMemory_9_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_9_fields_0 <= _GEN_3012;
          end
        end else if (_T_221) begin
          if (4'h9 == idxUpdate_6[3:0]) begin
            TBEMemory_9_fields_0 <= 32'h0;
          end else begin
            TBEMemory_9_fields_0 <= _GEN_3012;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'h9 == idxUpdate_6[3:0]) begin
              TBEMemory_9_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_9_fields_0 <= _GEN_3012;
            end
          end else begin
            TBEMemory_9_fields_0 <= _GEN_3012;
          end
        end else begin
          TBEMemory_9_fields_0 <= _GEN_3012;
        end
      end else if (isAlloc_6) begin
        if (4'h9 == idxAlloc[3:0]) begin
          TBEMemory_9_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_9_fields_0 <= _GEN_3012;
        end
      end else if (_T_221) begin
        if (4'h9 == idxUpdate_6[3:0]) begin
          TBEMemory_9_fields_0 <= 32'h0;
        end else begin
          TBEMemory_9_fields_0 <= _GEN_3012;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'h9 == idxUpdate_6[3:0]) begin
            TBEMemory_9_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_9_fields_0 <= _GEN_3012;
          end
        end else begin
          TBEMemory_9_fields_0 <= _GEN_3012;
        end
      end else begin
        TBEMemory_9_fields_0 <= _GEN_3012;
      end
    end else begin
      TBEMemory_9_fields_0 <= _GEN_3526;
    end
    if (reset) begin
      TBEMemory_10_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'ha == idxAlloc[3:0]) begin
        TBEMemory_10_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'ha == idxAlloc[3:0]) begin
          TBEMemory_10_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEMemory_10_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEMemory_10_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEMemory_10_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEMemory_10_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEMemory_10_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEMemory_10_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEMemory_10_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'ha == idxUpdate_0[3:0]) begin
                        TBEMemory_10_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEMemory_10_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEMemory_10_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'ha == idxUpdate_0[3:0]) begin
                        TBEMemory_10_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'ha == idxAlloc[3:0]) begin
                        TBEMemory_10_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'ha == idxUpdate_0[3:0]) begin
                        TBEMemory_10_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'ha == idxUpdate_0[3:0]) begin
                          TBEMemory_10_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEMemory_10_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEMemory_10_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'ha == idxUpdate_0[3:0]) begin
                        TBEMemory_10_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_10_state_state <= _GEN_475;
                end
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEMemory_10_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_10_state_state <= _GEN_475;
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_state_state <= 2'h0;
                  end else begin
                    TBEMemory_10_state_state <= _GEN_475;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_10_state_state <= _GEN_475;
                  end else if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_10_state_state <= _GEN_475;
                  end
                end else begin
                  TBEMemory_10_state_state <= _GEN_475;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEMemory_10_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_10_state_state <= _GEN_475;
                    end
                  end else if (_T_111) begin
                    if (4'ha == idxUpdate_1[3:0]) begin
                      TBEMemory_10_state_state <= 2'h0;
                    end else begin
                      TBEMemory_10_state_state <= _GEN_475;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_10_state_state <= _GEN_475;
                    end else if (4'ha == idxUpdate_1[3:0]) begin
                      TBEMemory_10_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_10_state_state <= _GEN_475;
                    end
                  end else begin
                    TBEMemory_10_state_state <= _GEN_475;
                  end
                end else if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEMemory_10_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_10_state_state <= _GEN_475;
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_state_state <= 2'h0;
                  end else begin
                    TBEMemory_10_state_state <= _GEN_475;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_10_state_state <= _GEN_475;
                  end else if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_10_state_state <= _GEN_475;
                  end
                end else begin
                  TBEMemory_10_state_state <= _GEN_475;
                end
              end else begin
                TBEMemory_10_state_state <= _GEN_989;
              end
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEMemory_10_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_10_state_state <= _GEN_989;
                end
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_state_state <= 2'h0;
                end else begin
                  TBEMemory_10_state_state <= _GEN_989;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_10_state_state <= _GEN_989;
                end else if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_10_state_state <= _GEN_989;
                end
              end else begin
                TBEMemory_10_state_state <= _GEN_989;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEMemory_10_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_10_state_state <= _GEN_989;
                  end
                end else if (_T_133) begin
                  if (4'ha == idxUpdate_2[3:0]) begin
                    TBEMemory_10_state_state <= 2'h0;
                  end else begin
                    TBEMemory_10_state_state <= _GEN_989;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_10_state_state <= _GEN_989;
                  end else if (4'ha == idxUpdate_2[3:0]) begin
                    TBEMemory_10_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_10_state_state <= _GEN_989;
                  end
                end else begin
                  TBEMemory_10_state_state <= _GEN_989;
                end
              end else if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEMemory_10_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_10_state_state <= _GEN_989;
                end
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_state_state <= 2'h0;
                end else begin
                  TBEMemory_10_state_state <= _GEN_989;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_10_state_state <= _GEN_989;
                end else if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_10_state_state <= _GEN_989;
                end
              end else begin
                TBEMemory_10_state_state <= _GEN_989;
              end
            end else begin
              TBEMemory_10_state_state <= _GEN_1503;
            end
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEMemory_10_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_10_state_state <= _GEN_1503;
              end
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_state_state <= 2'h0;
              end else begin
                TBEMemory_10_state_state <= _GEN_1503;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_10_state_state <= _GEN_1503;
              end else if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_10_state_state <= _GEN_1503;
              end
            end else begin
              TBEMemory_10_state_state <= _GEN_1503;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEMemory_10_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_10_state_state <= _GEN_1503;
                end
              end else if (_T_155) begin
                if (4'ha == idxUpdate_3[3:0]) begin
                  TBEMemory_10_state_state <= 2'h0;
                end else begin
                  TBEMemory_10_state_state <= _GEN_1503;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_10_state_state <= _GEN_1503;
                end else if (4'ha == idxUpdate_3[3:0]) begin
                  TBEMemory_10_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_10_state_state <= _GEN_1503;
                end
              end else begin
                TBEMemory_10_state_state <= _GEN_1503;
              end
            end else if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEMemory_10_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_10_state_state <= _GEN_1503;
              end
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_state_state <= 2'h0;
              end else begin
                TBEMemory_10_state_state <= _GEN_1503;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_10_state_state <= _GEN_1503;
              end else if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_10_state_state <= _GEN_1503;
              end
            end else begin
              TBEMemory_10_state_state <= _GEN_1503;
            end
          end else begin
            TBEMemory_10_state_state <= _GEN_2017;
          end
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEMemory_10_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_10_state_state <= _GEN_2017;
            end
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_state_state <= 2'h0;
            end else begin
              TBEMemory_10_state_state <= _GEN_2017;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_10_state_state <= _GEN_2017;
            end else if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_10_state_state <= _GEN_2017;
            end
          end else begin
            TBEMemory_10_state_state <= _GEN_2017;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEMemory_10_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_10_state_state <= _GEN_2017;
              end
            end else if (_T_177) begin
              if (4'ha == idxUpdate_4[3:0]) begin
                TBEMemory_10_state_state <= 2'h0;
              end else begin
                TBEMemory_10_state_state <= _GEN_2017;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_10_state_state <= _GEN_2017;
              end else if (4'ha == idxUpdate_4[3:0]) begin
                TBEMemory_10_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_10_state_state <= _GEN_2017;
              end
            end else begin
              TBEMemory_10_state_state <= _GEN_2017;
            end
          end else if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEMemory_10_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_10_state_state <= _GEN_2017;
            end
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_state_state <= 2'h0;
            end else begin
              TBEMemory_10_state_state <= _GEN_2017;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_10_state_state <= _GEN_2017;
            end else if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_10_state_state <= _GEN_2017;
            end
          end else begin
            TBEMemory_10_state_state <= _GEN_2017;
          end
        end else begin
          TBEMemory_10_state_state <= _GEN_2531;
        end
      end else if (_T_221) begin
        if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEMemory_10_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_10_state_state <= _GEN_2531;
          end
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_state_state <= 2'h0;
          end else begin
            TBEMemory_10_state_state <= _GEN_2531;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_10_state_state <= _GEN_2531;
          end else if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_10_state_state <= _GEN_2531;
          end
        end else begin
          TBEMemory_10_state_state <= _GEN_2531;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEMemory_10_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_10_state_state <= _GEN_2531;
            end
          end else if (_T_199) begin
            if (4'ha == idxUpdate_5[3:0]) begin
              TBEMemory_10_state_state <= 2'h0;
            end else begin
              TBEMemory_10_state_state <= _GEN_2531;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_10_state_state <= _GEN_2531;
            end else if (4'ha == idxUpdate_5[3:0]) begin
              TBEMemory_10_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_10_state_state <= _GEN_2531;
            end
          end else begin
            TBEMemory_10_state_state <= _GEN_2531;
          end
        end else if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEMemory_10_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_10_state_state <= _GEN_2531;
          end
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_state_state <= 2'h0;
          end else begin
            TBEMemory_10_state_state <= _GEN_2531;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_10_state_state <= _GEN_2531;
          end else if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_10_state_state <= _GEN_2531;
          end
        end else begin
          TBEMemory_10_state_state <= _GEN_2531;
        end
      end else begin
        TBEMemory_10_state_state <= _GEN_3045;
      end
    end else if (_T_243) begin
      if (4'ha == idxUpdate_7[3:0]) begin
        TBEMemory_10_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'ha == idxAlloc[3:0]) begin
          TBEMemory_10_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_10_state_state <= _GEN_3045;
        end
      end else if (_T_221) begin
        if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_state_state <= 2'h0;
        end else begin
          TBEMemory_10_state_state <= _GEN_3045;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_10_state_state <= _GEN_3045;
        end else if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_10_state_state <= _GEN_3045;
        end
      end else begin
        TBEMemory_10_state_state <= _GEN_3045;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEMemory_10_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_10_state_state <= _GEN_3045;
          end
        end else if (_T_221) begin
          if (4'ha == idxUpdate_6[3:0]) begin
            TBEMemory_10_state_state <= 2'h0;
          end else begin
            TBEMemory_10_state_state <= _GEN_3045;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_10_state_state <= _GEN_3045;
          end else if (4'ha == idxUpdate_6[3:0]) begin
            TBEMemory_10_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_10_state_state <= _GEN_3045;
          end
        end else begin
          TBEMemory_10_state_state <= _GEN_3045;
        end
      end else if (4'ha == idxUpdate_7[3:0]) begin
        TBEMemory_10_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'ha == idxAlloc[3:0]) begin
          TBEMemory_10_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_10_state_state <= _GEN_3045;
        end
      end else if (_T_221) begin
        if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_state_state <= 2'h0;
        end else begin
          TBEMemory_10_state_state <= _GEN_3045;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_10_state_state <= _GEN_3045;
        end else if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_10_state_state <= _GEN_3045;
        end
      end else begin
        TBEMemory_10_state_state <= _GEN_3045;
      end
    end else begin
      TBEMemory_10_state_state <= _GEN_3559;
    end
    if (reset) begin
      TBEMemory_10_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'ha == idxAlloc[3:0]) begin
        TBEMemory_10_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'ha == idxAlloc[3:0]) begin
          TBEMemory_10_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEMemory_10_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEMemory_10_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEMemory_10_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEMemory_10_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEMemory_10_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEMemory_10_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEMemory_10_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'ha == idxUpdate_0[3:0]) begin
                        TBEMemory_10_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEMemory_10_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEMemory_10_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'ha == idxUpdate_0[3:0]) begin
                        TBEMemory_10_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'ha == idxAlloc[3:0]) begin
                        TBEMemory_10_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'ha == idxUpdate_0[3:0]) begin
                        TBEMemory_10_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'ha == idxUpdate_0[3:0]) begin
                          TBEMemory_10_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEMemory_10_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEMemory_10_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'ha == idxUpdate_0[3:0]) begin
                        TBEMemory_10_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_10_way <= _GEN_459;
                end
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEMemory_10_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_10_way <= _GEN_459;
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_way <= 3'h2;
                  end else begin
                    TBEMemory_10_way <= _GEN_459;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_10_way <= _GEN_459;
                  end else if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_10_way <= _GEN_459;
                  end
                end else begin
                  TBEMemory_10_way <= _GEN_459;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEMemory_10_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_10_way <= _GEN_459;
                    end
                  end else if (_T_111) begin
                    if (4'ha == idxUpdate_1[3:0]) begin
                      TBEMemory_10_way <= 3'h2;
                    end else begin
                      TBEMemory_10_way <= _GEN_459;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_10_way <= _GEN_459;
                    end else if (4'ha == idxUpdate_1[3:0]) begin
                      TBEMemory_10_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_10_way <= _GEN_459;
                    end
                  end else begin
                    TBEMemory_10_way <= _GEN_459;
                  end
                end else if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEMemory_10_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_10_way <= _GEN_459;
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_way <= 3'h2;
                  end else begin
                    TBEMemory_10_way <= _GEN_459;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_10_way <= _GEN_459;
                  end else if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_10_way <= _GEN_459;
                  end
                end else begin
                  TBEMemory_10_way <= _GEN_459;
                end
              end else begin
                TBEMemory_10_way <= _GEN_973;
              end
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEMemory_10_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_10_way <= _GEN_973;
                end
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_way <= 3'h2;
                end else begin
                  TBEMemory_10_way <= _GEN_973;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_10_way <= _GEN_973;
                end else if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_10_way <= _GEN_973;
                end
              end else begin
                TBEMemory_10_way <= _GEN_973;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEMemory_10_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_10_way <= _GEN_973;
                  end
                end else if (_T_133) begin
                  if (4'ha == idxUpdate_2[3:0]) begin
                    TBEMemory_10_way <= 3'h2;
                  end else begin
                    TBEMemory_10_way <= _GEN_973;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_10_way <= _GEN_973;
                  end else if (4'ha == idxUpdate_2[3:0]) begin
                    TBEMemory_10_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_10_way <= _GEN_973;
                  end
                end else begin
                  TBEMemory_10_way <= _GEN_973;
                end
              end else if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEMemory_10_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_10_way <= _GEN_973;
                end
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_way <= 3'h2;
                end else begin
                  TBEMemory_10_way <= _GEN_973;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_10_way <= _GEN_973;
                end else if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_10_way <= _GEN_973;
                end
              end else begin
                TBEMemory_10_way <= _GEN_973;
              end
            end else begin
              TBEMemory_10_way <= _GEN_1487;
            end
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEMemory_10_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_10_way <= _GEN_1487;
              end
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_way <= 3'h2;
              end else begin
                TBEMemory_10_way <= _GEN_1487;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_10_way <= _GEN_1487;
              end else if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_10_way <= _GEN_1487;
              end
            end else begin
              TBEMemory_10_way <= _GEN_1487;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEMemory_10_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_10_way <= _GEN_1487;
                end
              end else if (_T_155) begin
                if (4'ha == idxUpdate_3[3:0]) begin
                  TBEMemory_10_way <= 3'h2;
                end else begin
                  TBEMemory_10_way <= _GEN_1487;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_10_way <= _GEN_1487;
                end else if (4'ha == idxUpdate_3[3:0]) begin
                  TBEMemory_10_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_10_way <= _GEN_1487;
                end
              end else begin
                TBEMemory_10_way <= _GEN_1487;
              end
            end else if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEMemory_10_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_10_way <= _GEN_1487;
              end
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_way <= 3'h2;
              end else begin
                TBEMemory_10_way <= _GEN_1487;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_10_way <= _GEN_1487;
              end else if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_10_way <= _GEN_1487;
              end
            end else begin
              TBEMemory_10_way <= _GEN_1487;
            end
          end else begin
            TBEMemory_10_way <= _GEN_2001;
          end
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEMemory_10_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_10_way <= _GEN_2001;
            end
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_way <= 3'h2;
            end else begin
              TBEMemory_10_way <= _GEN_2001;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_10_way <= _GEN_2001;
            end else if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_10_way <= _GEN_2001;
            end
          end else begin
            TBEMemory_10_way <= _GEN_2001;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEMemory_10_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_10_way <= _GEN_2001;
              end
            end else if (_T_177) begin
              if (4'ha == idxUpdate_4[3:0]) begin
                TBEMemory_10_way <= 3'h2;
              end else begin
                TBEMemory_10_way <= _GEN_2001;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_10_way <= _GEN_2001;
              end else if (4'ha == idxUpdate_4[3:0]) begin
                TBEMemory_10_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_10_way <= _GEN_2001;
              end
            end else begin
              TBEMemory_10_way <= _GEN_2001;
            end
          end else if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEMemory_10_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_10_way <= _GEN_2001;
            end
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_way <= 3'h2;
            end else begin
              TBEMemory_10_way <= _GEN_2001;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_10_way <= _GEN_2001;
            end else if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_10_way <= _GEN_2001;
            end
          end else begin
            TBEMemory_10_way <= _GEN_2001;
          end
        end else begin
          TBEMemory_10_way <= _GEN_2515;
        end
      end else if (_T_221) begin
        if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEMemory_10_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_10_way <= _GEN_2515;
          end
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_way <= 3'h2;
          end else begin
            TBEMemory_10_way <= _GEN_2515;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_10_way <= _GEN_2515;
          end else if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_10_way <= _GEN_2515;
          end
        end else begin
          TBEMemory_10_way <= _GEN_2515;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEMemory_10_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_10_way <= _GEN_2515;
            end
          end else if (_T_199) begin
            if (4'ha == idxUpdate_5[3:0]) begin
              TBEMemory_10_way <= 3'h2;
            end else begin
              TBEMemory_10_way <= _GEN_2515;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_10_way <= _GEN_2515;
            end else if (4'ha == idxUpdate_5[3:0]) begin
              TBEMemory_10_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_10_way <= _GEN_2515;
            end
          end else begin
            TBEMemory_10_way <= _GEN_2515;
          end
        end else if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEMemory_10_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_10_way <= _GEN_2515;
          end
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_way <= 3'h2;
          end else begin
            TBEMemory_10_way <= _GEN_2515;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_10_way <= _GEN_2515;
          end else if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_10_way <= _GEN_2515;
          end
        end else begin
          TBEMemory_10_way <= _GEN_2515;
        end
      end else begin
        TBEMemory_10_way <= _GEN_3029;
      end
    end else if (_T_243) begin
      if (4'ha == idxUpdate_7[3:0]) begin
        TBEMemory_10_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'ha == idxAlloc[3:0]) begin
          TBEMemory_10_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_10_way <= _GEN_3029;
        end
      end else if (_T_221) begin
        if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_way <= 3'h2;
        end else begin
          TBEMemory_10_way <= _GEN_3029;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_10_way <= _GEN_3029;
        end else if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_10_way <= _GEN_3029;
        end
      end else begin
        TBEMemory_10_way <= _GEN_3029;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEMemory_10_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_10_way <= _GEN_3029;
          end
        end else if (_T_221) begin
          if (4'ha == idxUpdate_6[3:0]) begin
            TBEMemory_10_way <= 3'h2;
          end else begin
            TBEMemory_10_way <= _GEN_3029;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_10_way <= _GEN_3029;
          end else if (4'ha == idxUpdate_6[3:0]) begin
            TBEMemory_10_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_10_way <= _GEN_3029;
          end
        end else begin
          TBEMemory_10_way <= _GEN_3029;
        end
      end else if (4'ha == idxUpdate_7[3:0]) begin
        TBEMemory_10_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'ha == idxAlloc[3:0]) begin
          TBEMemory_10_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_10_way <= _GEN_3029;
        end
      end else if (_T_221) begin
        if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_way <= 3'h2;
        end else begin
          TBEMemory_10_way <= _GEN_3029;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_10_way <= _GEN_3029;
        end else if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_10_way <= _GEN_3029;
        end
      end else begin
        TBEMemory_10_way <= _GEN_3029;
      end
    end else begin
      TBEMemory_10_way <= _GEN_3543;
    end
    if (reset) begin
      TBEMemory_10_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'ha == idxAlloc[3:0]) begin
        TBEMemory_10_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'ha == idxAlloc[3:0]) begin
          TBEMemory_10_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEMemory_10_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEMemory_10_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEMemory_10_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEMemory_10_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEMemory_10_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEMemory_10_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEMemory_10_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'ha == idxUpdate_0[3:0]) begin
                        TBEMemory_10_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEMemory_10_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEMemory_10_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'ha == idxUpdate_0[3:0]) begin
                        TBEMemory_10_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'ha == idxUpdate_1[3:0]) begin
                      TBEMemory_10_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'ha == idxAlloc[3:0]) begin
                        TBEMemory_10_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'ha == idxUpdate_0[3:0]) begin
                        TBEMemory_10_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'ha == idxUpdate_0[3:0]) begin
                          TBEMemory_10_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEMemory_10_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEMemory_10_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'ha == idxUpdate_0[3:0]) begin
                        TBEMemory_10_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_443;
                end
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEMemory_10_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_443;
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_443;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'ha == idxUpdate_1[3:0]) begin
                      TBEMemory_10_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_10_fields_0 <= _GEN_443;
                    end
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_443;
                  end
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_443;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'ha == idxUpdate_2[3:0]) begin
                    TBEMemory_10_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEMemory_10_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_10_fields_0 <= _GEN_443;
                    end
                  end else if (_T_111) begin
                    if (4'ha == idxUpdate_1[3:0]) begin
                      TBEMemory_10_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_10_fields_0 <= _GEN_443;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'ha == idxUpdate_1[3:0]) begin
                        TBEMemory_10_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_10_fields_0 <= _GEN_443;
                      end
                    end else begin
                      TBEMemory_10_fields_0 <= _GEN_443;
                    end
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_443;
                  end
                end else if (isAlloc_1) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEMemory_10_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_443;
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEMemory_10_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_443;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'ha == idxUpdate_1[3:0]) begin
                      TBEMemory_10_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_10_fields_0 <= _GEN_443;
                    end
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_443;
                  end
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_443;
                end
              end else begin
                TBEMemory_10_fields_0 <= _GEN_957;
              end
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEMemory_10_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_957;
                end
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_957;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'ha == idxUpdate_2[3:0]) begin
                    TBEMemory_10_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_957;
                  end
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_957;
                end
              end else begin
                TBEMemory_10_fields_0 <= _GEN_957;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'ha == idxUpdate_3[3:0]) begin
                  TBEMemory_10_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEMemory_10_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_957;
                  end
                end else if (_T_133) begin
                  if (4'ha == idxUpdate_2[3:0]) begin
                    TBEMemory_10_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_957;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'ha == idxUpdate_2[3:0]) begin
                      TBEMemory_10_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_10_fields_0 <= _GEN_957;
                    end
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_957;
                  end
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_957;
                end
              end else if (isAlloc_2) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEMemory_10_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_957;
                end
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEMemory_10_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_957;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'ha == idxUpdate_2[3:0]) begin
                    TBEMemory_10_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_957;
                  end
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_957;
                end
              end else begin
                TBEMemory_10_fields_0 <= _GEN_957;
              end
            end else begin
              TBEMemory_10_fields_0 <= _GEN_1471;
            end
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEMemory_10_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_10_fields_0 <= _GEN_1471;
              end
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_fields_0 <= 32'h0;
              end else begin
                TBEMemory_10_fields_0 <= _GEN_1471;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'ha == idxUpdate_3[3:0]) begin
                  TBEMemory_10_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_1471;
                end
              end else begin
                TBEMemory_10_fields_0 <= _GEN_1471;
              end
            end else begin
              TBEMemory_10_fields_0 <= _GEN_1471;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'ha == idxUpdate_4[3:0]) begin
                TBEMemory_10_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEMemory_10_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_1471;
                end
              end else if (_T_155) begin
                if (4'ha == idxUpdate_3[3:0]) begin
                  TBEMemory_10_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_1471;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'ha == idxUpdate_3[3:0]) begin
                    TBEMemory_10_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_10_fields_0 <= _GEN_1471;
                  end
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_1471;
                end
              end else begin
                TBEMemory_10_fields_0 <= _GEN_1471;
              end
            end else if (isAlloc_3) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEMemory_10_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_10_fields_0 <= _GEN_1471;
              end
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEMemory_10_fields_0 <= 32'h0;
              end else begin
                TBEMemory_10_fields_0 <= _GEN_1471;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'ha == idxUpdate_3[3:0]) begin
                  TBEMemory_10_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_1471;
                end
              end else begin
                TBEMemory_10_fields_0 <= _GEN_1471;
              end
            end else begin
              TBEMemory_10_fields_0 <= _GEN_1471;
            end
          end else begin
            TBEMemory_10_fields_0 <= _GEN_1985;
          end
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEMemory_10_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_10_fields_0 <= _GEN_1985;
            end
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_fields_0 <= 32'h0;
            end else begin
              TBEMemory_10_fields_0 <= _GEN_1985;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'ha == idxUpdate_4[3:0]) begin
                TBEMemory_10_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_10_fields_0 <= _GEN_1985;
              end
            end else begin
              TBEMemory_10_fields_0 <= _GEN_1985;
            end
          end else begin
            TBEMemory_10_fields_0 <= _GEN_1985;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'ha == idxUpdate_5[3:0]) begin
              TBEMemory_10_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEMemory_10_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_10_fields_0 <= _GEN_1985;
              end
            end else if (_T_177) begin
              if (4'ha == idxUpdate_4[3:0]) begin
                TBEMemory_10_fields_0 <= 32'h0;
              end else begin
                TBEMemory_10_fields_0 <= _GEN_1985;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'ha == idxUpdate_4[3:0]) begin
                  TBEMemory_10_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_10_fields_0 <= _GEN_1985;
                end
              end else begin
                TBEMemory_10_fields_0 <= _GEN_1985;
              end
            end else begin
              TBEMemory_10_fields_0 <= _GEN_1985;
            end
          end else if (isAlloc_4) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEMemory_10_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_10_fields_0 <= _GEN_1985;
            end
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEMemory_10_fields_0 <= 32'h0;
            end else begin
              TBEMemory_10_fields_0 <= _GEN_1985;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'ha == idxUpdate_4[3:0]) begin
                TBEMemory_10_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_10_fields_0 <= _GEN_1985;
              end
            end else begin
              TBEMemory_10_fields_0 <= _GEN_1985;
            end
          end else begin
            TBEMemory_10_fields_0 <= _GEN_1985;
          end
        end else begin
          TBEMemory_10_fields_0 <= _GEN_2499;
        end
      end else if (_T_221) begin
        if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEMemory_10_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_10_fields_0 <= _GEN_2499;
          end
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_fields_0 <= 32'h0;
          end else begin
            TBEMemory_10_fields_0 <= _GEN_2499;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'ha == idxUpdate_5[3:0]) begin
              TBEMemory_10_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_10_fields_0 <= _GEN_2499;
            end
          end else begin
            TBEMemory_10_fields_0 <= _GEN_2499;
          end
        end else begin
          TBEMemory_10_fields_0 <= _GEN_2499;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'ha == idxUpdate_6[3:0]) begin
            TBEMemory_10_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEMemory_10_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_10_fields_0 <= _GEN_2499;
            end
          end else if (_T_199) begin
            if (4'ha == idxUpdate_5[3:0]) begin
              TBEMemory_10_fields_0 <= 32'h0;
            end else begin
              TBEMemory_10_fields_0 <= _GEN_2499;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'ha == idxUpdate_5[3:0]) begin
                TBEMemory_10_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_10_fields_0 <= _GEN_2499;
              end
            end else begin
              TBEMemory_10_fields_0 <= _GEN_2499;
            end
          end else begin
            TBEMemory_10_fields_0 <= _GEN_2499;
          end
        end else if (isAlloc_5) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEMemory_10_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_10_fields_0 <= _GEN_2499;
          end
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEMemory_10_fields_0 <= 32'h0;
          end else begin
            TBEMemory_10_fields_0 <= _GEN_2499;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'ha == idxUpdate_5[3:0]) begin
              TBEMemory_10_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_10_fields_0 <= _GEN_2499;
            end
          end else begin
            TBEMemory_10_fields_0 <= _GEN_2499;
          end
        end else begin
          TBEMemory_10_fields_0 <= _GEN_2499;
        end
      end else begin
        TBEMemory_10_fields_0 <= _GEN_3013;
      end
    end else if (_T_243) begin
      if (4'ha == idxUpdate_7[3:0]) begin
        TBEMemory_10_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'ha == idxAlloc[3:0]) begin
          TBEMemory_10_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_10_fields_0 <= _GEN_3013;
        end
      end else if (_T_221) begin
        if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_fields_0 <= 32'h0;
        end else begin
          TBEMemory_10_fields_0 <= _GEN_3013;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'ha == idxUpdate_6[3:0]) begin
            TBEMemory_10_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_10_fields_0 <= _GEN_3013;
          end
        end else begin
          TBEMemory_10_fields_0 <= _GEN_3013;
        end
      end else begin
        TBEMemory_10_fields_0 <= _GEN_3013;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'ha == idxUpdate_7[3:0]) begin
          TBEMemory_10_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEMemory_10_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_10_fields_0 <= _GEN_3013;
          end
        end else if (_T_221) begin
          if (4'ha == idxUpdate_6[3:0]) begin
            TBEMemory_10_fields_0 <= 32'h0;
          end else begin
            TBEMemory_10_fields_0 <= _GEN_3013;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'ha == idxUpdate_6[3:0]) begin
              TBEMemory_10_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_10_fields_0 <= _GEN_3013;
            end
          end else begin
            TBEMemory_10_fields_0 <= _GEN_3013;
          end
        end else begin
          TBEMemory_10_fields_0 <= _GEN_3013;
        end
      end else if (isAlloc_6) begin
        if (4'ha == idxAlloc[3:0]) begin
          TBEMemory_10_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_10_fields_0 <= _GEN_3013;
        end
      end else if (_T_221) begin
        if (4'ha == idxUpdate_6[3:0]) begin
          TBEMemory_10_fields_0 <= 32'h0;
        end else begin
          TBEMemory_10_fields_0 <= _GEN_3013;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'ha == idxUpdate_6[3:0]) begin
            TBEMemory_10_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_10_fields_0 <= _GEN_3013;
          end
        end else begin
          TBEMemory_10_fields_0 <= _GEN_3013;
        end
      end else begin
        TBEMemory_10_fields_0 <= _GEN_3013;
      end
    end else begin
      TBEMemory_10_fields_0 <= _GEN_3527;
    end
    if (reset) begin
      TBEMemory_11_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'hb == idxAlloc[3:0]) begin
        TBEMemory_11_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'hb == idxAlloc[3:0]) begin
          TBEMemory_11_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEMemory_11_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEMemory_11_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEMemory_11_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEMemory_11_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEMemory_11_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEMemory_11_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEMemory_11_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hb == idxUpdate_0[3:0]) begin
                        TBEMemory_11_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEMemory_11_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEMemory_11_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hb == idxUpdate_0[3:0]) begin
                        TBEMemory_11_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'hb == idxAlloc[3:0]) begin
                        TBEMemory_11_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'hb == idxUpdate_0[3:0]) begin
                        TBEMemory_11_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'hb == idxUpdate_0[3:0]) begin
                          TBEMemory_11_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEMemory_11_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEMemory_11_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hb == idxUpdate_0[3:0]) begin
                        TBEMemory_11_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_11_state_state <= _GEN_476;
                end
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEMemory_11_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_11_state_state <= _GEN_476;
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_state_state <= 2'h0;
                  end else begin
                    TBEMemory_11_state_state <= _GEN_476;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_11_state_state <= _GEN_476;
                  end else if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_11_state_state <= _GEN_476;
                  end
                end else begin
                  TBEMemory_11_state_state <= _GEN_476;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEMemory_11_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_11_state_state <= _GEN_476;
                    end
                  end else if (_T_111) begin
                    if (4'hb == idxUpdate_1[3:0]) begin
                      TBEMemory_11_state_state <= 2'h0;
                    end else begin
                      TBEMemory_11_state_state <= _GEN_476;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_11_state_state <= _GEN_476;
                    end else if (4'hb == idxUpdate_1[3:0]) begin
                      TBEMemory_11_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_11_state_state <= _GEN_476;
                    end
                  end else begin
                    TBEMemory_11_state_state <= _GEN_476;
                  end
                end else if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEMemory_11_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_11_state_state <= _GEN_476;
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_state_state <= 2'h0;
                  end else begin
                    TBEMemory_11_state_state <= _GEN_476;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_11_state_state <= _GEN_476;
                  end else if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_11_state_state <= _GEN_476;
                  end
                end else begin
                  TBEMemory_11_state_state <= _GEN_476;
                end
              end else begin
                TBEMemory_11_state_state <= _GEN_990;
              end
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEMemory_11_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_11_state_state <= _GEN_990;
                end
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_state_state <= 2'h0;
                end else begin
                  TBEMemory_11_state_state <= _GEN_990;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_11_state_state <= _GEN_990;
                end else if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_11_state_state <= _GEN_990;
                end
              end else begin
                TBEMemory_11_state_state <= _GEN_990;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEMemory_11_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_11_state_state <= _GEN_990;
                  end
                end else if (_T_133) begin
                  if (4'hb == idxUpdate_2[3:0]) begin
                    TBEMemory_11_state_state <= 2'h0;
                  end else begin
                    TBEMemory_11_state_state <= _GEN_990;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_11_state_state <= _GEN_990;
                  end else if (4'hb == idxUpdate_2[3:0]) begin
                    TBEMemory_11_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_11_state_state <= _GEN_990;
                  end
                end else begin
                  TBEMemory_11_state_state <= _GEN_990;
                end
              end else if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEMemory_11_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_11_state_state <= _GEN_990;
                end
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_state_state <= 2'h0;
                end else begin
                  TBEMemory_11_state_state <= _GEN_990;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_11_state_state <= _GEN_990;
                end else if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_11_state_state <= _GEN_990;
                end
              end else begin
                TBEMemory_11_state_state <= _GEN_990;
              end
            end else begin
              TBEMemory_11_state_state <= _GEN_1504;
            end
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEMemory_11_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_11_state_state <= _GEN_1504;
              end
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_state_state <= 2'h0;
              end else begin
                TBEMemory_11_state_state <= _GEN_1504;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_11_state_state <= _GEN_1504;
              end else if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_11_state_state <= _GEN_1504;
              end
            end else begin
              TBEMemory_11_state_state <= _GEN_1504;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEMemory_11_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_11_state_state <= _GEN_1504;
                end
              end else if (_T_155) begin
                if (4'hb == idxUpdate_3[3:0]) begin
                  TBEMemory_11_state_state <= 2'h0;
                end else begin
                  TBEMemory_11_state_state <= _GEN_1504;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_11_state_state <= _GEN_1504;
                end else if (4'hb == idxUpdate_3[3:0]) begin
                  TBEMemory_11_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_11_state_state <= _GEN_1504;
                end
              end else begin
                TBEMemory_11_state_state <= _GEN_1504;
              end
            end else if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEMemory_11_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_11_state_state <= _GEN_1504;
              end
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_state_state <= 2'h0;
              end else begin
                TBEMemory_11_state_state <= _GEN_1504;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_11_state_state <= _GEN_1504;
              end else if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_11_state_state <= _GEN_1504;
              end
            end else begin
              TBEMemory_11_state_state <= _GEN_1504;
            end
          end else begin
            TBEMemory_11_state_state <= _GEN_2018;
          end
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEMemory_11_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_11_state_state <= _GEN_2018;
            end
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_state_state <= 2'h0;
            end else begin
              TBEMemory_11_state_state <= _GEN_2018;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_11_state_state <= _GEN_2018;
            end else if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_11_state_state <= _GEN_2018;
            end
          end else begin
            TBEMemory_11_state_state <= _GEN_2018;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEMemory_11_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_11_state_state <= _GEN_2018;
              end
            end else if (_T_177) begin
              if (4'hb == idxUpdate_4[3:0]) begin
                TBEMemory_11_state_state <= 2'h0;
              end else begin
                TBEMemory_11_state_state <= _GEN_2018;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_11_state_state <= _GEN_2018;
              end else if (4'hb == idxUpdate_4[3:0]) begin
                TBEMemory_11_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_11_state_state <= _GEN_2018;
              end
            end else begin
              TBEMemory_11_state_state <= _GEN_2018;
            end
          end else if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEMemory_11_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_11_state_state <= _GEN_2018;
            end
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_state_state <= 2'h0;
            end else begin
              TBEMemory_11_state_state <= _GEN_2018;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_11_state_state <= _GEN_2018;
            end else if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_11_state_state <= _GEN_2018;
            end
          end else begin
            TBEMemory_11_state_state <= _GEN_2018;
          end
        end else begin
          TBEMemory_11_state_state <= _GEN_2532;
        end
      end else if (_T_221) begin
        if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEMemory_11_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_11_state_state <= _GEN_2532;
          end
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_state_state <= 2'h0;
          end else begin
            TBEMemory_11_state_state <= _GEN_2532;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_11_state_state <= _GEN_2532;
          end else if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_11_state_state <= _GEN_2532;
          end
        end else begin
          TBEMemory_11_state_state <= _GEN_2532;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEMemory_11_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_11_state_state <= _GEN_2532;
            end
          end else if (_T_199) begin
            if (4'hb == idxUpdate_5[3:0]) begin
              TBEMemory_11_state_state <= 2'h0;
            end else begin
              TBEMemory_11_state_state <= _GEN_2532;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_11_state_state <= _GEN_2532;
            end else if (4'hb == idxUpdate_5[3:0]) begin
              TBEMemory_11_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_11_state_state <= _GEN_2532;
            end
          end else begin
            TBEMemory_11_state_state <= _GEN_2532;
          end
        end else if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEMemory_11_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_11_state_state <= _GEN_2532;
          end
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_state_state <= 2'h0;
          end else begin
            TBEMemory_11_state_state <= _GEN_2532;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_11_state_state <= _GEN_2532;
          end else if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_11_state_state <= _GEN_2532;
          end
        end else begin
          TBEMemory_11_state_state <= _GEN_2532;
        end
      end else begin
        TBEMemory_11_state_state <= _GEN_3046;
      end
    end else if (_T_243) begin
      if (4'hb == idxUpdate_7[3:0]) begin
        TBEMemory_11_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'hb == idxAlloc[3:0]) begin
          TBEMemory_11_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_11_state_state <= _GEN_3046;
        end
      end else if (_T_221) begin
        if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_state_state <= 2'h0;
        end else begin
          TBEMemory_11_state_state <= _GEN_3046;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_11_state_state <= _GEN_3046;
        end else if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_11_state_state <= _GEN_3046;
        end
      end else begin
        TBEMemory_11_state_state <= _GEN_3046;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEMemory_11_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_11_state_state <= _GEN_3046;
          end
        end else if (_T_221) begin
          if (4'hb == idxUpdate_6[3:0]) begin
            TBEMemory_11_state_state <= 2'h0;
          end else begin
            TBEMemory_11_state_state <= _GEN_3046;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_11_state_state <= _GEN_3046;
          end else if (4'hb == idxUpdate_6[3:0]) begin
            TBEMemory_11_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_11_state_state <= _GEN_3046;
          end
        end else begin
          TBEMemory_11_state_state <= _GEN_3046;
        end
      end else if (4'hb == idxUpdate_7[3:0]) begin
        TBEMemory_11_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'hb == idxAlloc[3:0]) begin
          TBEMemory_11_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_11_state_state <= _GEN_3046;
        end
      end else if (_T_221) begin
        if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_state_state <= 2'h0;
        end else begin
          TBEMemory_11_state_state <= _GEN_3046;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_11_state_state <= _GEN_3046;
        end else if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_11_state_state <= _GEN_3046;
        end
      end else begin
        TBEMemory_11_state_state <= _GEN_3046;
      end
    end else begin
      TBEMemory_11_state_state <= _GEN_3560;
    end
    if (reset) begin
      TBEMemory_11_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'hb == idxAlloc[3:0]) begin
        TBEMemory_11_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'hb == idxAlloc[3:0]) begin
          TBEMemory_11_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEMemory_11_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEMemory_11_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEMemory_11_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEMemory_11_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEMemory_11_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEMemory_11_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEMemory_11_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hb == idxUpdate_0[3:0]) begin
                        TBEMemory_11_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEMemory_11_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEMemory_11_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hb == idxUpdate_0[3:0]) begin
                        TBEMemory_11_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'hb == idxAlloc[3:0]) begin
                        TBEMemory_11_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'hb == idxUpdate_0[3:0]) begin
                        TBEMemory_11_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'hb == idxUpdate_0[3:0]) begin
                          TBEMemory_11_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEMemory_11_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEMemory_11_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hb == idxUpdate_0[3:0]) begin
                        TBEMemory_11_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_11_way <= _GEN_460;
                end
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEMemory_11_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_11_way <= _GEN_460;
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_way <= 3'h2;
                  end else begin
                    TBEMemory_11_way <= _GEN_460;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_11_way <= _GEN_460;
                  end else if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_11_way <= _GEN_460;
                  end
                end else begin
                  TBEMemory_11_way <= _GEN_460;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEMemory_11_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_11_way <= _GEN_460;
                    end
                  end else if (_T_111) begin
                    if (4'hb == idxUpdate_1[3:0]) begin
                      TBEMemory_11_way <= 3'h2;
                    end else begin
                      TBEMemory_11_way <= _GEN_460;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_11_way <= _GEN_460;
                    end else if (4'hb == idxUpdate_1[3:0]) begin
                      TBEMemory_11_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_11_way <= _GEN_460;
                    end
                  end else begin
                    TBEMemory_11_way <= _GEN_460;
                  end
                end else if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEMemory_11_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_11_way <= _GEN_460;
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_way <= 3'h2;
                  end else begin
                    TBEMemory_11_way <= _GEN_460;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_11_way <= _GEN_460;
                  end else if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_11_way <= _GEN_460;
                  end
                end else begin
                  TBEMemory_11_way <= _GEN_460;
                end
              end else begin
                TBEMemory_11_way <= _GEN_974;
              end
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEMemory_11_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_11_way <= _GEN_974;
                end
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_way <= 3'h2;
                end else begin
                  TBEMemory_11_way <= _GEN_974;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_11_way <= _GEN_974;
                end else if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_11_way <= _GEN_974;
                end
              end else begin
                TBEMemory_11_way <= _GEN_974;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEMemory_11_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_11_way <= _GEN_974;
                  end
                end else if (_T_133) begin
                  if (4'hb == idxUpdate_2[3:0]) begin
                    TBEMemory_11_way <= 3'h2;
                  end else begin
                    TBEMemory_11_way <= _GEN_974;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_11_way <= _GEN_974;
                  end else if (4'hb == idxUpdate_2[3:0]) begin
                    TBEMemory_11_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_11_way <= _GEN_974;
                  end
                end else begin
                  TBEMemory_11_way <= _GEN_974;
                end
              end else if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEMemory_11_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_11_way <= _GEN_974;
                end
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_way <= 3'h2;
                end else begin
                  TBEMemory_11_way <= _GEN_974;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_11_way <= _GEN_974;
                end else if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_11_way <= _GEN_974;
                end
              end else begin
                TBEMemory_11_way <= _GEN_974;
              end
            end else begin
              TBEMemory_11_way <= _GEN_1488;
            end
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEMemory_11_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_11_way <= _GEN_1488;
              end
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_way <= 3'h2;
              end else begin
                TBEMemory_11_way <= _GEN_1488;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_11_way <= _GEN_1488;
              end else if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_11_way <= _GEN_1488;
              end
            end else begin
              TBEMemory_11_way <= _GEN_1488;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEMemory_11_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_11_way <= _GEN_1488;
                end
              end else if (_T_155) begin
                if (4'hb == idxUpdate_3[3:0]) begin
                  TBEMemory_11_way <= 3'h2;
                end else begin
                  TBEMemory_11_way <= _GEN_1488;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_11_way <= _GEN_1488;
                end else if (4'hb == idxUpdate_3[3:0]) begin
                  TBEMemory_11_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_11_way <= _GEN_1488;
                end
              end else begin
                TBEMemory_11_way <= _GEN_1488;
              end
            end else if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEMemory_11_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_11_way <= _GEN_1488;
              end
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_way <= 3'h2;
              end else begin
                TBEMemory_11_way <= _GEN_1488;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_11_way <= _GEN_1488;
              end else if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_11_way <= _GEN_1488;
              end
            end else begin
              TBEMemory_11_way <= _GEN_1488;
            end
          end else begin
            TBEMemory_11_way <= _GEN_2002;
          end
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEMemory_11_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_11_way <= _GEN_2002;
            end
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_way <= 3'h2;
            end else begin
              TBEMemory_11_way <= _GEN_2002;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_11_way <= _GEN_2002;
            end else if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_11_way <= _GEN_2002;
            end
          end else begin
            TBEMemory_11_way <= _GEN_2002;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEMemory_11_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_11_way <= _GEN_2002;
              end
            end else if (_T_177) begin
              if (4'hb == idxUpdate_4[3:0]) begin
                TBEMemory_11_way <= 3'h2;
              end else begin
                TBEMemory_11_way <= _GEN_2002;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_11_way <= _GEN_2002;
              end else if (4'hb == idxUpdate_4[3:0]) begin
                TBEMemory_11_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_11_way <= _GEN_2002;
              end
            end else begin
              TBEMemory_11_way <= _GEN_2002;
            end
          end else if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEMemory_11_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_11_way <= _GEN_2002;
            end
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_way <= 3'h2;
            end else begin
              TBEMemory_11_way <= _GEN_2002;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_11_way <= _GEN_2002;
            end else if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_11_way <= _GEN_2002;
            end
          end else begin
            TBEMemory_11_way <= _GEN_2002;
          end
        end else begin
          TBEMemory_11_way <= _GEN_2516;
        end
      end else if (_T_221) begin
        if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEMemory_11_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_11_way <= _GEN_2516;
          end
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_way <= 3'h2;
          end else begin
            TBEMemory_11_way <= _GEN_2516;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_11_way <= _GEN_2516;
          end else if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_11_way <= _GEN_2516;
          end
        end else begin
          TBEMemory_11_way <= _GEN_2516;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEMemory_11_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_11_way <= _GEN_2516;
            end
          end else if (_T_199) begin
            if (4'hb == idxUpdate_5[3:0]) begin
              TBEMemory_11_way <= 3'h2;
            end else begin
              TBEMemory_11_way <= _GEN_2516;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_11_way <= _GEN_2516;
            end else if (4'hb == idxUpdate_5[3:0]) begin
              TBEMemory_11_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_11_way <= _GEN_2516;
            end
          end else begin
            TBEMemory_11_way <= _GEN_2516;
          end
        end else if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEMemory_11_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_11_way <= _GEN_2516;
          end
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_way <= 3'h2;
          end else begin
            TBEMemory_11_way <= _GEN_2516;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_11_way <= _GEN_2516;
          end else if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_11_way <= _GEN_2516;
          end
        end else begin
          TBEMemory_11_way <= _GEN_2516;
        end
      end else begin
        TBEMemory_11_way <= _GEN_3030;
      end
    end else if (_T_243) begin
      if (4'hb == idxUpdate_7[3:0]) begin
        TBEMemory_11_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'hb == idxAlloc[3:0]) begin
          TBEMemory_11_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_11_way <= _GEN_3030;
        end
      end else if (_T_221) begin
        if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_way <= 3'h2;
        end else begin
          TBEMemory_11_way <= _GEN_3030;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_11_way <= _GEN_3030;
        end else if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_11_way <= _GEN_3030;
        end
      end else begin
        TBEMemory_11_way <= _GEN_3030;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEMemory_11_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_11_way <= _GEN_3030;
          end
        end else if (_T_221) begin
          if (4'hb == idxUpdate_6[3:0]) begin
            TBEMemory_11_way <= 3'h2;
          end else begin
            TBEMemory_11_way <= _GEN_3030;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_11_way <= _GEN_3030;
          end else if (4'hb == idxUpdate_6[3:0]) begin
            TBEMemory_11_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_11_way <= _GEN_3030;
          end
        end else begin
          TBEMemory_11_way <= _GEN_3030;
        end
      end else if (4'hb == idxUpdate_7[3:0]) begin
        TBEMemory_11_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'hb == idxAlloc[3:0]) begin
          TBEMemory_11_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_11_way <= _GEN_3030;
        end
      end else if (_T_221) begin
        if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_way <= 3'h2;
        end else begin
          TBEMemory_11_way <= _GEN_3030;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_11_way <= _GEN_3030;
        end else if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_11_way <= _GEN_3030;
        end
      end else begin
        TBEMemory_11_way <= _GEN_3030;
      end
    end else begin
      TBEMemory_11_way <= _GEN_3544;
    end
    if (reset) begin
      TBEMemory_11_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'hb == idxAlloc[3:0]) begin
        TBEMemory_11_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'hb == idxAlloc[3:0]) begin
          TBEMemory_11_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEMemory_11_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEMemory_11_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEMemory_11_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEMemory_11_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEMemory_11_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEMemory_11_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEMemory_11_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'hb == idxUpdate_0[3:0]) begin
                        TBEMemory_11_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEMemory_11_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEMemory_11_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'hb == idxUpdate_0[3:0]) begin
                        TBEMemory_11_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'hb == idxUpdate_1[3:0]) begin
                      TBEMemory_11_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'hb == idxAlloc[3:0]) begin
                        TBEMemory_11_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'hb == idxUpdate_0[3:0]) begin
                        TBEMemory_11_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'hb == idxUpdate_0[3:0]) begin
                          TBEMemory_11_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEMemory_11_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEMemory_11_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'hb == idxUpdate_0[3:0]) begin
                        TBEMemory_11_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_444;
                end
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEMemory_11_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_444;
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_444;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'hb == idxUpdate_1[3:0]) begin
                      TBEMemory_11_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_11_fields_0 <= _GEN_444;
                    end
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_444;
                  end
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_444;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'hb == idxUpdate_2[3:0]) begin
                    TBEMemory_11_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEMemory_11_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_11_fields_0 <= _GEN_444;
                    end
                  end else if (_T_111) begin
                    if (4'hb == idxUpdate_1[3:0]) begin
                      TBEMemory_11_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_11_fields_0 <= _GEN_444;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'hb == idxUpdate_1[3:0]) begin
                        TBEMemory_11_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_11_fields_0 <= _GEN_444;
                      end
                    end else begin
                      TBEMemory_11_fields_0 <= _GEN_444;
                    end
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_444;
                  end
                end else if (isAlloc_1) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEMemory_11_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_444;
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEMemory_11_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_444;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'hb == idxUpdate_1[3:0]) begin
                      TBEMemory_11_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_11_fields_0 <= _GEN_444;
                    end
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_444;
                  end
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_444;
                end
              end else begin
                TBEMemory_11_fields_0 <= _GEN_958;
              end
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEMemory_11_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_958;
                end
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_958;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'hb == idxUpdate_2[3:0]) begin
                    TBEMemory_11_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_958;
                  end
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_958;
                end
              end else begin
                TBEMemory_11_fields_0 <= _GEN_958;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'hb == idxUpdate_3[3:0]) begin
                  TBEMemory_11_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEMemory_11_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_958;
                  end
                end else if (_T_133) begin
                  if (4'hb == idxUpdate_2[3:0]) begin
                    TBEMemory_11_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_958;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'hb == idxUpdate_2[3:0]) begin
                      TBEMemory_11_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_11_fields_0 <= _GEN_958;
                    end
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_958;
                  end
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_958;
                end
              end else if (isAlloc_2) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEMemory_11_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_958;
                end
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEMemory_11_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_958;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'hb == idxUpdate_2[3:0]) begin
                    TBEMemory_11_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_958;
                  end
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_958;
                end
              end else begin
                TBEMemory_11_fields_0 <= _GEN_958;
              end
            end else begin
              TBEMemory_11_fields_0 <= _GEN_1472;
            end
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEMemory_11_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_11_fields_0 <= _GEN_1472;
              end
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_fields_0 <= 32'h0;
              end else begin
                TBEMemory_11_fields_0 <= _GEN_1472;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'hb == idxUpdate_3[3:0]) begin
                  TBEMemory_11_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_1472;
                end
              end else begin
                TBEMemory_11_fields_0 <= _GEN_1472;
              end
            end else begin
              TBEMemory_11_fields_0 <= _GEN_1472;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'hb == idxUpdate_4[3:0]) begin
                TBEMemory_11_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEMemory_11_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_1472;
                end
              end else if (_T_155) begin
                if (4'hb == idxUpdate_3[3:0]) begin
                  TBEMemory_11_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_1472;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'hb == idxUpdate_3[3:0]) begin
                    TBEMemory_11_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_11_fields_0 <= _GEN_1472;
                  end
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_1472;
                end
              end else begin
                TBEMemory_11_fields_0 <= _GEN_1472;
              end
            end else if (isAlloc_3) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEMemory_11_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_11_fields_0 <= _GEN_1472;
              end
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEMemory_11_fields_0 <= 32'h0;
              end else begin
                TBEMemory_11_fields_0 <= _GEN_1472;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'hb == idxUpdate_3[3:0]) begin
                  TBEMemory_11_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_1472;
                end
              end else begin
                TBEMemory_11_fields_0 <= _GEN_1472;
              end
            end else begin
              TBEMemory_11_fields_0 <= _GEN_1472;
            end
          end else begin
            TBEMemory_11_fields_0 <= _GEN_1986;
          end
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEMemory_11_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_11_fields_0 <= _GEN_1986;
            end
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_fields_0 <= 32'h0;
            end else begin
              TBEMemory_11_fields_0 <= _GEN_1986;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'hb == idxUpdate_4[3:0]) begin
                TBEMemory_11_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_11_fields_0 <= _GEN_1986;
              end
            end else begin
              TBEMemory_11_fields_0 <= _GEN_1986;
            end
          end else begin
            TBEMemory_11_fields_0 <= _GEN_1986;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'hb == idxUpdate_5[3:0]) begin
              TBEMemory_11_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEMemory_11_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_11_fields_0 <= _GEN_1986;
              end
            end else if (_T_177) begin
              if (4'hb == idxUpdate_4[3:0]) begin
                TBEMemory_11_fields_0 <= 32'h0;
              end else begin
                TBEMemory_11_fields_0 <= _GEN_1986;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'hb == idxUpdate_4[3:0]) begin
                  TBEMemory_11_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_11_fields_0 <= _GEN_1986;
                end
              end else begin
                TBEMemory_11_fields_0 <= _GEN_1986;
              end
            end else begin
              TBEMemory_11_fields_0 <= _GEN_1986;
            end
          end else if (isAlloc_4) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEMemory_11_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_11_fields_0 <= _GEN_1986;
            end
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEMemory_11_fields_0 <= 32'h0;
            end else begin
              TBEMemory_11_fields_0 <= _GEN_1986;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'hb == idxUpdate_4[3:0]) begin
                TBEMemory_11_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_11_fields_0 <= _GEN_1986;
              end
            end else begin
              TBEMemory_11_fields_0 <= _GEN_1986;
            end
          end else begin
            TBEMemory_11_fields_0 <= _GEN_1986;
          end
        end else begin
          TBEMemory_11_fields_0 <= _GEN_2500;
        end
      end else if (_T_221) begin
        if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEMemory_11_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_11_fields_0 <= _GEN_2500;
          end
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_fields_0 <= 32'h0;
          end else begin
            TBEMemory_11_fields_0 <= _GEN_2500;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'hb == idxUpdate_5[3:0]) begin
              TBEMemory_11_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_11_fields_0 <= _GEN_2500;
            end
          end else begin
            TBEMemory_11_fields_0 <= _GEN_2500;
          end
        end else begin
          TBEMemory_11_fields_0 <= _GEN_2500;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'hb == idxUpdate_6[3:0]) begin
            TBEMemory_11_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEMemory_11_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_11_fields_0 <= _GEN_2500;
            end
          end else if (_T_199) begin
            if (4'hb == idxUpdate_5[3:0]) begin
              TBEMemory_11_fields_0 <= 32'h0;
            end else begin
              TBEMemory_11_fields_0 <= _GEN_2500;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'hb == idxUpdate_5[3:0]) begin
                TBEMemory_11_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_11_fields_0 <= _GEN_2500;
              end
            end else begin
              TBEMemory_11_fields_0 <= _GEN_2500;
            end
          end else begin
            TBEMemory_11_fields_0 <= _GEN_2500;
          end
        end else if (isAlloc_5) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEMemory_11_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_11_fields_0 <= _GEN_2500;
          end
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEMemory_11_fields_0 <= 32'h0;
          end else begin
            TBEMemory_11_fields_0 <= _GEN_2500;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'hb == idxUpdate_5[3:0]) begin
              TBEMemory_11_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_11_fields_0 <= _GEN_2500;
            end
          end else begin
            TBEMemory_11_fields_0 <= _GEN_2500;
          end
        end else begin
          TBEMemory_11_fields_0 <= _GEN_2500;
        end
      end else begin
        TBEMemory_11_fields_0 <= _GEN_3014;
      end
    end else if (_T_243) begin
      if (4'hb == idxUpdate_7[3:0]) begin
        TBEMemory_11_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'hb == idxAlloc[3:0]) begin
          TBEMemory_11_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_11_fields_0 <= _GEN_3014;
        end
      end else if (_T_221) begin
        if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_fields_0 <= 32'h0;
        end else begin
          TBEMemory_11_fields_0 <= _GEN_3014;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'hb == idxUpdate_6[3:0]) begin
            TBEMemory_11_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_11_fields_0 <= _GEN_3014;
          end
        end else begin
          TBEMemory_11_fields_0 <= _GEN_3014;
        end
      end else begin
        TBEMemory_11_fields_0 <= _GEN_3014;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'hb == idxUpdate_7[3:0]) begin
          TBEMemory_11_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEMemory_11_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_11_fields_0 <= _GEN_3014;
          end
        end else if (_T_221) begin
          if (4'hb == idxUpdate_6[3:0]) begin
            TBEMemory_11_fields_0 <= 32'h0;
          end else begin
            TBEMemory_11_fields_0 <= _GEN_3014;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'hb == idxUpdate_6[3:0]) begin
              TBEMemory_11_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_11_fields_0 <= _GEN_3014;
            end
          end else begin
            TBEMemory_11_fields_0 <= _GEN_3014;
          end
        end else begin
          TBEMemory_11_fields_0 <= _GEN_3014;
        end
      end else if (isAlloc_6) begin
        if (4'hb == idxAlloc[3:0]) begin
          TBEMemory_11_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_11_fields_0 <= _GEN_3014;
        end
      end else if (_T_221) begin
        if (4'hb == idxUpdate_6[3:0]) begin
          TBEMemory_11_fields_0 <= 32'h0;
        end else begin
          TBEMemory_11_fields_0 <= _GEN_3014;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'hb == idxUpdate_6[3:0]) begin
            TBEMemory_11_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_11_fields_0 <= _GEN_3014;
          end
        end else begin
          TBEMemory_11_fields_0 <= _GEN_3014;
        end
      end else begin
        TBEMemory_11_fields_0 <= _GEN_3014;
      end
    end else begin
      TBEMemory_11_fields_0 <= _GEN_3528;
    end
    if (reset) begin
      TBEMemory_12_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'hc == idxAlloc[3:0]) begin
        TBEMemory_12_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'hc == idxAlloc[3:0]) begin
          TBEMemory_12_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEMemory_12_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEMemory_12_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEMemory_12_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEMemory_12_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEMemory_12_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEMemory_12_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEMemory_12_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hc == idxUpdate_0[3:0]) begin
                        TBEMemory_12_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEMemory_12_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEMemory_12_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hc == idxUpdate_0[3:0]) begin
                        TBEMemory_12_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'hc == idxAlloc[3:0]) begin
                        TBEMemory_12_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'hc == idxUpdate_0[3:0]) begin
                        TBEMemory_12_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'hc == idxUpdate_0[3:0]) begin
                          TBEMemory_12_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEMemory_12_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEMemory_12_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hc == idxUpdate_0[3:0]) begin
                        TBEMemory_12_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_12_state_state <= _GEN_477;
                end
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEMemory_12_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_12_state_state <= _GEN_477;
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_state_state <= 2'h0;
                  end else begin
                    TBEMemory_12_state_state <= _GEN_477;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_12_state_state <= _GEN_477;
                  end else if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_12_state_state <= _GEN_477;
                  end
                end else begin
                  TBEMemory_12_state_state <= _GEN_477;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEMemory_12_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_12_state_state <= _GEN_477;
                    end
                  end else if (_T_111) begin
                    if (4'hc == idxUpdate_1[3:0]) begin
                      TBEMemory_12_state_state <= 2'h0;
                    end else begin
                      TBEMemory_12_state_state <= _GEN_477;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_12_state_state <= _GEN_477;
                    end else if (4'hc == idxUpdate_1[3:0]) begin
                      TBEMemory_12_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_12_state_state <= _GEN_477;
                    end
                  end else begin
                    TBEMemory_12_state_state <= _GEN_477;
                  end
                end else if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEMemory_12_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_12_state_state <= _GEN_477;
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_state_state <= 2'h0;
                  end else begin
                    TBEMemory_12_state_state <= _GEN_477;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_12_state_state <= _GEN_477;
                  end else if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_12_state_state <= _GEN_477;
                  end
                end else begin
                  TBEMemory_12_state_state <= _GEN_477;
                end
              end else begin
                TBEMemory_12_state_state <= _GEN_991;
              end
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEMemory_12_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_12_state_state <= _GEN_991;
                end
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_state_state <= 2'h0;
                end else begin
                  TBEMemory_12_state_state <= _GEN_991;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_12_state_state <= _GEN_991;
                end else if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_12_state_state <= _GEN_991;
                end
              end else begin
                TBEMemory_12_state_state <= _GEN_991;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEMemory_12_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_12_state_state <= _GEN_991;
                  end
                end else if (_T_133) begin
                  if (4'hc == idxUpdate_2[3:0]) begin
                    TBEMemory_12_state_state <= 2'h0;
                  end else begin
                    TBEMemory_12_state_state <= _GEN_991;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_12_state_state <= _GEN_991;
                  end else if (4'hc == idxUpdate_2[3:0]) begin
                    TBEMemory_12_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_12_state_state <= _GEN_991;
                  end
                end else begin
                  TBEMemory_12_state_state <= _GEN_991;
                end
              end else if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEMemory_12_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_12_state_state <= _GEN_991;
                end
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_state_state <= 2'h0;
                end else begin
                  TBEMemory_12_state_state <= _GEN_991;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_12_state_state <= _GEN_991;
                end else if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_12_state_state <= _GEN_991;
                end
              end else begin
                TBEMemory_12_state_state <= _GEN_991;
              end
            end else begin
              TBEMemory_12_state_state <= _GEN_1505;
            end
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEMemory_12_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_12_state_state <= _GEN_1505;
              end
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_state_state <= 2'h0;
              end else begin
                TBEMemory_12_state_state <= _GEN_1505;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_12_state_state <= _GEN_1505;
              end else if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_12_state_state <= _GEN_1505;
              end
            end else begin
              TBEMemory_12_state_state <= _GEN_1505;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEMemory_12_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_12_state_state <= _GEN_1505;
                end
              end else if (_T_155) begin
                if (4'hc == idxUpdate_3[3:0]) begin
                  TBEMemory_12_state_state <= 2'h0;
                end else begin
                  TBEMemory_12_state_state <= _GEN_1505;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_12_state_state <= _GEN_1505;
                end else if (4'hc == idxUpdate_3[3:0]) begin
                  TBEMemory_12_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_12_state_state <= _GEN_1505;
                end
              end else begin
                TBEMemory_12_state_state <= _GEN_1505;
              end
            end else if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEMemory_12_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_12_state_state <= _GEN_1505;
              end
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_state_state <= 2'h0;
              end else begin
                TBEMemory_12_state_state <= _GEN_1505;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_12_state_state <= _GEN_1505;
              end else if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_12_state_state <= _GEN_1505;
              end
            end else begin
              TBEMemory_12_state_state <= _GEN_1505;
            end
          end else begin
            TBEMemory_12_state_state <= _GEN_2019;
          end
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEMemory_12_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_12_state_state <= _GEN_2019;
            end
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_state_state <= 2'h0;
            end else begin
              TBEMemory_12_state_state <= _GEN_2019;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_12_state_state <= _GEN_2019;
            end else if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_12_state_state <= _GEN_2019;
            end
          end else begin
            TBEMemory_12_state_state <= _GEN_2019;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEMemory_12_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_12_state_state <= _GEN_2019;
              end
            end else if (_T_177) begin
              if (4'hc == idxUpdate_4[3:0]) begin
                TBEMemory_12_state_state <= 2'h0;
              end else begin
                TBEMemory_12_state_state <= _GEN_2019;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_12_state_state <= _GEN_2019;
              end else if (4'hc == idxUpdate_4[3:0]) begin
                TBEMemory_12_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_12_state_state <= _GEN_2019;
              end
            end else begin
              TBEMemory_12_state_state <= _GEN_2019;
            end
          end else if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEMemory_12_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_12_state_state <= _GEN_2019;
            end
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_state_state <= 2'h0;
            end else begin
              TBEMemory_12_state_state <= _GEN_2019;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_12_state_state <= _GEN_2019;
            end else if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_12_state_state <= _GEN_2019;
            end
          end else begin
            TBEMemory_12_state_state <= _GEN_2019;
          end
        end else begin
          TBEMemory_12_state_state <= _GEN_2533;
        end
      end else if (_T_221) begin
        if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEMemory_12_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_12_state_state <= _GEN_2533;
          end
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_state_state <= 2'h0;
          end else begin
            TBEMemory_12_state_state <= _GEN_2533;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_12_state_state <= _GEN_2533;
          end else if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_12_state_state <= _GEN_2533;
          end
        end else begin
          TBEMemory_12_state_state <= _GEN_2533;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEMemory_12_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_12_state_state <= _GEN_2533;
            end
          end else if (_T_199) begin
            if (4'hc == idxUpdate_5[3:0]) begin
              TBEMemory_12_state_state <= 2'h0;
            end else begin
              TBEMemory_12_state_state <= _GEN_2533;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_12_state_state <= _GEN_2533;
            end else if (4'hc == idxUpdate_5[3:0]) begin
              TBEMemory_12_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_12_state_state <= _GEN_2533;
            end
          end else begin
            TBEMemory_12_state_state <= _GEN_2533;
          end
        end else if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEMemory_12_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_12_state_state <= _GEN_2533;
          end
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_state_state <= 2'h0;
          end else begin
            TBEMemory_12_state_state <= _GEN_2533;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_12_state_state <= _GEN_2533;
          end else if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_12_state_state <= _GEN_2533;
          end
        end else begin
          TBEMemory_12_state_state <= _GEN_2533;
        end
      end else begin
        TBEMemory_12_state_state <= _GEN_3047;
      end
    end else if (_T_243) begin
      if (4'hc == idxUpdate_7[3:0]) begin
        TBEMemory_12_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'hc == idxAlloc[3:0]) begin
          TBEMemory_12_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_12_state_state <= _GEN_3047;
        end
      end else if (_T_221) begin
        if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_state_state <= 2'h0;
        end else begin
          TBEMemory_12_state_state <= _GEN_3047;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_12_state_state <= _GEN_3047;
        end else if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_12_state_state <= _GEN_3047;
        end
      end else begin
        TBEMemory_12_state_state <= _GEN_3047;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEMemory_12_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_12_state_state <= _GEN_3047;
          end
        end else if (_T_221) begin
          if (4'hc == idxUpdate_6[3:0]) begin
            TBEMemory_12_state_state <= 2'h0;
          end else begin
            TBEMemory_12_state_state <= _GEN_3047;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_12_state_state <= _GEN_3047;
          end else if (4'hc == idxUpdate_6[3:0]) begin
            TBEMemory_12_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_12_state_state <= _GEN_3047;
          end
        end else begin
          TBEMemory_12_state_state <= _GEN_3047;
        end
      end else if (4'hc == idxUpdate_7[3:0]) begin
        TBEMemory_12_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'hc == idxAlloc[3:0]) begin
          TBEMemory_12_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_12_state_state <= _GEN_3047;
        end
      end else if (_T_221) begin
        if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_state_state <= 2'h0;
        end else begin
          TBEMemory_12_state_state <= _GEN_3047;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_12_state_state <= _GEN_3047;
        end else if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_12_state_state <= _GEN_3047;
        end
      end else begin
        TBEMemory_12_state_state <= _GEN_3047;
      end
    end else begin
      TBEMemory_12_state_state <= _GEN_3561;
    end
    if (reset) begin
      TBEMemory_12_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'hc == idxAlloc[3:0]) begin
        TBEMemory_12_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'hc == idxAlloc[3:0]) begin
          TBEMemory_12_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEMemory_12_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEMemory_12_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEMemory_12_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEMemory_12_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEMemory_12_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEMemory_12_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEMemory_12_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hc == idxUpdate_0[3:0]) begin
                        TBEMemory_12_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEMemory_12_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEMemory_12_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hc == idxUpdate_0[3:0]) begin
                        TBEMemory_12_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'hc == idxAlloc[3:0]) begin
                        TBEMemory_12_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'hc == idxUpdate_0[3:0]) begin
                        TBEMemory_12_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'hc == idxUpdate_0[3:0]) begin
                          TBEMemory_12_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEMemory_12_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEMemory_12_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hc == idxUpdate_0[3:0]) begin
                        TBEMemory_12_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_12_way <= _GEN_461;
                end
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEMemory_12_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_12_way <= _GEN_461;
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_way <= 3'h2;
                  end else begin
                    TBEMemory_12_way <= _GEN_461;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_12_way <= _GEN_461;
                  end else if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_12_way <= _GEN_461;
                  end
                end else begin
                  TBEMemory_12_way <= _GEN_461;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEMemory_12_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_12_way <= _GEN_461;
                    end
                  end else if (_T_111) begin
                    if (4'hc == idxUpdate_1[3:0]) begin
                      TBEMemory_12_way <= 3'h2;
                    end else begin
                      TBEMemory_12_way <= _GEN_461;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_12_way <= _GEN_461;
                    end else if (4'hc == idxUpdate_1[3:0]) begin
                      TBEMemory_12_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_12_way <= _GEN_461;
                    end
                  end else begin
                    TBEMemory_12_way <= _GEN_461;
                  end
                end else if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEMemory_12_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_12_way <= _GEN_461;
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_way <= 3'h2;
                  end else begin
                    TBEMemory_12_way <= _GEN_461;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_12_way <= _GEN_461;
                  end else if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_12_way <= _GEN_461;
                  end
                end else begin
                  TBEMemory_12_way <= _GEN_461;
                end
              end else begin
                TBEMemory_12_way <= _GEN_975;
              end
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEMemory_12_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_12_way <= _GEN_975;
                end
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_way <= 3'h2;
                end else begin
                  TBEMemory_12_way <= _GEN_975;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_12_way <= _GEN_975;
                end else if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_12_way <= _GEN_975;
                end
              end else begin
                TBEMemory_12_way <= _GEN_975;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEMemory_12_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_12_way <= _GEN_975;
                  end
                end else if (_T_133) begin
                  if (4'hc == idxUpdate_2[3:0]) begin
                    TBEMemory_12_way <= 3'h2;
                  end else begin
                    TBEMemory_12_way <= _GEN_975;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_12_way <= _GEN_975;
                  end else if (4'hc == idxUpdate_2[3:0]) begin
                    TBEMemory_12_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_12_way <= _GEN_975;
                  end
                end else begin
                  TBEMemory_12_way <= _GEN_975;
                end
              end else if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEMemory_12_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_12_way <= _GEN_975;
                end
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_way <= 3'h2;
                end else begin
                  TBEMemory_12_way <= _GEN_975;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_12_way <= _GEN_975;
                end else if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_12_way <= _GEN_975;
                end
              end else begin
                TBEMemory_12_way <= _GEN_975;
              end
            end else begin
              TBEMemory_12_way <= _GEN_1489;
            end
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEMemory_12_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_12_way <= _GEN_1489;
              end
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_way <= 3'h2;
              end else begin
                TBEMemory_12_way <= _GEN_1489;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_12_way <= _GEN_1489;
              end else if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_12_way <= _GEN_1489;
              end
            end else begin
              TBEMemory_12_way <= _GEN_1489;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEMemory_12_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_12_way <= _GEN_1489;
                end
              end else if (_T_155) begin
                if (4'hc == idxUpdate_3[3:0]) begin
                  TBEMemory_12_way <= 3'h2;
                end else begin
                  TBEMemory_12_way <= _GEN_1489;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_12_way <= _GEN_1489;
                end else if (4'hc == idxUpdate_3[3:0]) begin
                  TBEMemory_12_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_12_way <= _GEN_1489;
                end
              end else begin
                TBEMemory_12_way <= _GEN_1489;
              end
            end else if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEMemory_12_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_12_way <= _GEN_1489;
              end
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_way <= 3'h2;
              end else begin
                TBEMemory_12_way <= _GEN_1489;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_12_way <= _GEN_1489;
              end else if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_12_way <= _GEN_1489;
              end
            end else begin
              TBEMemory_12_way <= _GEN_1489;
            end
          end else begin
            TBEMemory_12_way <= _GEN_2003;
          end
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEMemory_12_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_12_way <= _GEN_2003;
            end
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_way <= 3'h2;
            end else begin
              TBEMemory_12_way <= _GEN_2003;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_12_way <= _GEN_2003;
            end else if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_12_way <= _GEN_2003;
            end
          end else begin
            TBEMemory_12_way <= _GEN_2003;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEMemory_12_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_12_way <= _GEN_2003;
              end
            end else if (_T_177) begin
              if (4'hc == idxUpdate_4[3:0]) begin
                TBEMemory_12_way <= 3'h2;
              end else begin
                TBEMemory_12_way <= _GEN_2003;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_12_way <= _GEN_2003;
              end else if (4'hc == idxUpdate_4[3:0]) begin
                TBEMemory_12_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_12_way <= _GEN_2003;
              end
            end else begin
              TBEMemory_12_way <= _GEN_2003;
            end
          end else if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEMemory_12_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_12_way <= _GEN_2003;
            end
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_way <= 3'h2;
            end else begin
              TBEMemory_12_way <= _GEN_2003;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_12_way <= _GEN_2003;
            end else if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_12_way <= _GEN_2003;
            end
          end else begin
            TBEMemory_12_way <= _GEN_2003;
          end
        end else begin
          TBEMemory_12_way <= _GEN_2517;
        end
      end else if (_T_221) begin
        if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEMemory_12_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_12_way <= _GEN_2517;
          end
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_way <= 3'h2;
          end else begin
            TBEMemory_12_way <= _GEN_2517;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_12_way <= _GEN_2517;
          end else if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_12_way <= _GEN_2517;
          end
        end else begin
          TBEMemory_12_way <= _GEN_2517;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEMemory_12_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_12_way <= _GEN_2517;
            end
          end else if (_T_199) begin
            if (4'hc == idxUpdate_5[3:0]) begin
              TBEMemory_12_way <= 3'h2;
            end else begin
              TBEMemory_12_way <= _GEN_2517;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_12_way <= _GEN_2517;
            end else if (4'hc == idxUpdate_5[3:0]) begin
              TBEMemory_12_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_12_way <= _GEN_2517;
            end
          end else begin
            TBEMemory_12_way <= _GEN_2517;
          end
        end else if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEMemory_12_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_12_way <= _GEN_2517;
          end
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_way <= 3'h2;
          end else begin
            TBEMemory_12_way <= _GEN_2517;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_12_way <= _GEN_2517;
          end else if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_12_way <= _GEN_2517;
          end
        end else begin
          TBEMemory_12_way <= _GEN_2517;
        end
      end else begin
        TBEMemory_12_way <= _GEN_3031;
      end
    end else if (_T_243) begin
      if (4'hc == idxUpdate_7[3:0]) begin
        TBEMemory_12_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'hc == idxAlloc[3:0]) begin
          TBEMemory_12_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_12_way <= _GEN_3031;
        end
      end else if (_T_221) begin
        if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_way <= 3'h2;
        end else begin
          TBEMemory_12_way <= _GEN_3031;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_12_way <= _GEN_3031;
        end else if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_12_way <= _GEN_3031;
        end
      end else begin
        TBEMemory_12_way <= _GEN_3031;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEMemory_12_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_12_way <= _GEN_3031;
          end
        end else if (_T_221) begin
          if (4'hc == idxUpdate_6[3:0]) begin
            TBEMemory_12_way <= 3'h2;
          end else begin
            TBEMemory_12_way <= _GEN_3031;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_12_way <= _GEN_3031;
          end else if (4'hc == idxUpdate_6[3:0]) begin
            TBEMemory_12_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_12_way <= _GEN_3031;
          end
        end else begin
          TBEMemory_12_way <= _GEN_3031;
        end
      end else if (4'hc == idxUpdate_7[3:0]) begin
        TBEMemory_12_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'hc == idxAlloc[3:0]) begin
          TBEMemory_12_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_12_way <= _GEN_3031;
        end
      end else if (_T_221) begin
        if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_way <= 3'h2;
        end else begin
          TBEMemory_12_way <= _GEN_3031;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_12_way <= _GEN_3031;
        end else if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_12_way <= _GEN_3031;
        end
      end else begin
        TBEMemory_12_way <= _GEN_3031;
      end
    end else begin
      TBEMemory_12_way <= _GEN_3545;
    end
    if (reset) begin
      TBEMemory_12_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'hc == idxAlloc[3:0]) begin
        TBEMemory_12_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'hc == idxAlloc[3:0]) begin
          TBEMemory_12_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEMemory_12_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEMemory_12_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEMemory_12_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEMemory_12_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEMemory_12_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEMemory_12_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEMemory_12_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'hc == idxUpdate_0[3:0]) begin
                        TBEMemory_12_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEMemory_12_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEMemory_12_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'hc == idxUpdate_0[3:0]) begin
                        TBEMemory_12_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'hc == idxUpdate_1[3:0]) begin
                      TBEMemory_12_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'hc == idxAlloc[3:0]) begin
                        TBEMemory_12_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'hc == idxUpdate_0[3:0]) begin
                        TBEMemory_12_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'hc == idxUpdate_0[3:0]) begin
                          TBEMemory_12_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEMemory_12_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEMemory_12_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'hc == idxUpdate_0[3:0]) begin
                        TBEMemory_12_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_445;
                end
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEMemory_12_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_445;
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_445;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'hc == idxUpdate_1[3:0]) begin
                      TBEMemory_12_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_12_fields_0 <= _GEN_445;
                    end
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_445;
                  end
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_445;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'hc == idxUpdate_2[3:0]) begin
                    TBEMemory_12_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEMemory_12_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_12_fields_0 <= _GEN_445;
                    end
                  end else if (_T_111) begin
                    if (4'hc == idxUpdate_1[3:0]) begin
                      TBEMemory_12_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_12_fields_0 <= _GEN_445;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'hc == idxUpdate_1[3:0]) begin
                        TBEMemory_12_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_12_fields_0 <= _GEN_445;
                      end
                    end else begin
                      TBEMemory_12_fields_0 <= _GEN_445;
                    end
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_445;
                  end
                end else if (isAlloc_1) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEMemory_12_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_445;
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEMemory_12_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_445;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'hc == idxUpdate_1[3:0]) begin
                      TBEMemory_12_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_12_fields_0 <= _GEN_445;
                    end
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_445;
                  end
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_445;
                end
              end else begin
                TBEMemory_12_fields_0 <= _GEN_959;
              end
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEMemory_12_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_959;
                end
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_959;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'hc == idxUpdate_2[3:0]) begin
                    TBEMemory_12_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_959;
                  end
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_959;
                end
              end else begin
                TBEMemory_12_fields_0 <= _GEN_959;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'hc == idxUpdate_3[3:0]) begin
                  TBEMemory_12_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEMemory_12_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_959;
                  end
                end else if (_T_133) begin
                  if (4'hc == idxUpdate_2[3:0]) begin
                    TBEMemory_12_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_959;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'hc == idxUpdate_2[3:0]) begin
                      TBEMemory_12_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_12_fields_0 <= _GEN_959;
                    end
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_959;
                  end
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_959;
                end
              end else if (isAlloc_2) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEMemory_12_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_959;
                end
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEMemory_12_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_959;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'hc == idxUpdate_2[3:0]) begin
                    TBEMemory_12_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_959;
                  end
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_959;
                end
              end else begin
                TBEMemory_12_fields_0 <= _GEN_959;
              end
            end else begin
              TBEMemory_12_fields_0 <= _GEN_1473;
            end
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEMemory_12_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_12_fields_0 <= _GEN_1473;
              end
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_fields_0 <= 32'h0;
              end else begin
                TBEMemory_12_fields_0 <= _GEN_1473;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'hc == idxUpdate_3[3:0]) begin
                  TBEMemory_12_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_1473;
                end
              end else begin
                TBEMemory_12_fields_0 <= _GEN_1473;
              end
            end else begin
              TBEMemory_12_fields_0 <= _GEN_1473;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'hc == idxUpdate_4[3:0]) begin
                TBEMemory_12_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEMemory_12_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_1473;
                end
              end else if (_T_155) begin
                if (4'hc == idxUpdate_3[3:0]) begin
                  TBEMemory_12_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_1473;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'hc == idxUpdate_3[3:0]) begin
                    TBEMemory_12_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_12_fields_0 <= _GEN_1473;
                  end
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_1473;
                end
              end else begin
                TBEMemory_12_fields_0 <= _GEN_1473;
              end
            end else if (isAlloc_3) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEMemory_12_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_12_fields_0 <= _GEN_1473;
              end
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEMemory_12_fields_0 <= 32'h0;
              end else begin
                TBEMemory_12_fields_0 <= _GEN_1473;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'hc == idxUpdate_3[3:0]) begin
                  TBEMemory_12_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_1473;
                end
              end else begin
                TBEMemory_12_fields_0 <= _GEN_1473;
              end
            end else begin
              TBEMemory_12_fields_0 <= _GEN_1473;
            end
          end else begin
            TBEMemory_12_fields_0 <= _GEN_1987;
          end
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEMemory_12_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_12_fields_0 <= _GEN_1987;
            end
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_fields_0 <= 32'h0;
            end else begin
              TBEMemory_12_fields_0 <= _GEN_1987;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'hc == idxUpdate_4[3:0]) begin
                TBEMemory_12_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_12_fields_0 <= _GEN_1987;
              end
            end else begin
              TBEMemory_12_fields_0 <= _GEN_1987;
            end
          end else begin
            TBEMemory_12_fields_0 <= _GEN_1987;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'hc == idxUpdate_5[3:0]) begin
              TBEMemory_12_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEMemory_12_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_12_fields_0 <= _GEN_1987;
              end
            end else if (_T_177) begin
              if (4'hc == idxUpdate_4[3:0]) begin
                TBEMemory_12_fields_0 <= 32'h0;
              end else begin
                TBEMemory_12_fields_0 <= _GEN_1987;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'hc == idxUpdate_4[3:0]) begin
                  TBEMemory_12_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_12_fields_0 <= _GEN_1987;
                end
              end else begin
                TBEMemory_12_fields_0 <= _GEN_1987;
              end
            end else begin
              TBEMemory_12_fields_0 <= _GEN_1987;
            end
          end else if (isAlloc_4) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEMemory_12_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_12_fields_0 <= _GEN_1987;
            end
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEMemory_12_fields_0 <= 32'h0;
            end else begin
              TBEMemory_12_fields_0 <= _GEN_1987;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'hc == idxUpdate_4[3:0]) begin
                TBEMemory_12_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_12_fields_0 <= _GEN_1987;
              end
            end else begin
              TBEMemory_12_fields_0 <= _GEN_1987;
            end
          end else begin
            TBEMemory_12_fields_0 <= _GEN_1987;
          end
        end else begin
          TBEMemory_12_fields_0 <= _GEN_2501;
        end
      end else if (_T_221) begin
        if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEMemory_12_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_12_fields_0 <= _GEN_2501;
          end
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_fields_0 <= 32'h0;
          end else begin
            TBEMemory_12_fields_0 <= _GEN_2501;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'hc == idxUpdate_5[3:0]) begin
              TBEMemory_12_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_12_fields_0 <= _GEN_2501;
            end
          end else begin
            TBEMemory_12_fields_0 <= _GEN_2501;
          end
        end else begin
          TBEMemory_12_fields_0 <= _GEN_2501;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'hc == idxUpdate_6[3:0]) begin
            TBEMemory_12_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEMemory_12_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_12_fields_0 <= _GEN_2501;
            end
          end else if (_T_199) begin
            if (4'hc == idxUpdate_5[3:0]) begin
              TBEMemory_12_fields_0 <= 32'h0;
            end else begin
              TBEMemory_12_fields_0 <= _GEN_2501;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'hc == idxUpdate_5[3:0]) begin
                TBEMemory_12_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_12_fields_0 <= _GEN_2501;
              end
            end else begin
              TBEMemory_12_fields_0 <= _GEN_2501;
            end
          end else begin
            TBEMemory_12_fields_0 <= _GEN_2501;
          end
        end else if (isAlloc_5) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEMemory_12_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_12_fields_0 <= _GEN_2501;
          end
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEMemory_12_fields_0 <= 32'h0;
          end else begin
            TBEMemory_12_fields_0 <= _GEN_2501;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'hc == idxUpdate_5[3:0]) begin
              TBEMemory_12_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_12_fields_0 <= _GEN_2501;
            end
          end else begin
            TBEMemory_12_fields_0 <= _GEN_2501;
          end
        end else begin
          TBEMemory_12_fields_0 <= _GEN_2501;
        end
      end else begin
        TBEMemory_12_fields_0 <= _GEN_3015;
      end
    end else if (_T_243) begin
      if (4'hc == idxUpdate_7[3:0]) begin
        TBEMemory_12_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'hc == idxAlloc[3:0]) begin
          TBEMemory_12_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_12_fields_0 <= _GEN_3015;
        end
      end else if (_T_221) begin
        if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_fields_0 <= 32'h0;
        end else begin
          TBEMemory_12_fields_0 <= _GEN_3015;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'hc == idxUpdate_6[3:0]) begin
            TBEMemory_12_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_12_fields_0 <= _GEN_3015;
          end
        end else begin
          TBEMemory_12_fields_0 <= _GEN_3015;
        end
      end else begin
        TBEMemory_12_fields_0 <= _GEN_3015;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'hc == idxUpdate_7[3:0]) begin
          TBEMemory_12_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEMemory_12_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_12_fields_0 <= _GEN_3015;
          end
        end else if (_T_221) begin
          if (4'hc == idxUpdate_6[3:0]) begin
            TBEMemory_12_fields_0 <= 32'h0;
          end else begin
            TBEMemory_12_fields_0 <= _GEN_3015;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'hc == idxUpdate_6[3:0]) begin
              TBEMemory_12_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_12_fields_0 <= _GEN_3015;
            end
          end else begin
            TBEMemory_12_fields_0 <= _GEN_3015;
          end
        end else begin
          TBEMemory_12_fields_0 <= _GEN_3015;
        end
      end else if (isAlloc_6) begin
        if (4'hc == idxAlloc[3:0]) begin
          TBEMemory_12_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_12_fields_0 <= _GEN_3015;
        end
      end else if (_T_221) begin
        if (4'hc == idxUpdate_6[3:0]) begin
          TBEMemory_12_fields_0 <= 32'h0;
        end else begin
          TBEMemory_12_fields_0 <= _GEN_3015;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'hc == idxUpdate_6[3:0]) begin
            TBEMemory_12_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_12_fields_0 <= _GEN_3015;
          end
        end else begin
          TBEMemory_12_fields_0 <= _GEN_3015;
        end
      end else begin
        TBEMemory_12_fields_0 <= _GEN_3015;
      end
    end else begin
      TBEMemory_12_fields_0 <= _GEN_3529;
    end
    if (reset) begin
      TBEMemory_13_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'hd == idxAlloc[3:0]) begin
        TBEMemory_13_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'hd == idxAlloc[3:0]) begin
          TBEMemory_13_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEMemory_13_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEMemory_13_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEMemory_13_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEMemory_13_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEMemory_13_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEMemory_13_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEMemory_13_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hd == idxUpdate_0[3:0]) begin
                        TBEMemory_13_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEMemory_13_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEMemory_13_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hd == idxUpdate_0[3:0]) begin
                        TBEMemory_13_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'hd == idxAlloc[3:0]) begin
                        TBEMemory_13_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'hd == idxUpdate_0[3:0]) begin
                        TBEMemory_13_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'hd == idxUpdate_0[3:0]) begin
                          TBEMemory_13_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEMemory_13_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEMemory_13_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hd == idxUpdate_0[3:0]) begin
                        TBEMemory_13_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_13_state_state <= _GEN_478;
                end
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEMemory_13_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_13_state_state <= _GEN_478;
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_state_state <= 2'h0;
                  end else begin
                    TBEMemory_13_state_state <= _GEN_478;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_13_state_state <= _GEN_478;
                  end else if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_13_state_state <= _GEN_478;
                  end
                end else begin
                  TBEMemory_13_state_state <= _GEN_478;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEMemory_13_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_13_state_state <= _GEN_478;
                    end
                  end else if (_T_111) begin
                    if (4'hd == idxUpdate_1[3:0]) begin
                      TBEMemory_13_state_state <= 2'h0;
                    end else begin
                      TBEMemory_13_state_state <= _GEN_478;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_13_state_state <= _GEN_478;
                    end else if (4'hd == idxUpdate_1[3:0]) begin
                      TBEMemory_13_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_13_state_state <= _GEN_478;
                    end
                  end else begin
                    TBEMemory_13_state_state <= _GEN_478;
                  end
                end else if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEMemory_13_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_13_state_state <= _GEN_478;
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_state_state <= 2'h0;
                  end else begin
                    TBEMemory_13_state_state <= _GEN_478;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_13_state_state <= _GEN_478;
                  end else if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_13_state_state <= _GEN_478;
                  end
                end else begin
                  TBEMemory_13_state_state <= _GEN_478;
                end
              end else begin
                TBEMemory_13_state_state <= _GEN_992;
              end
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEMemory_13_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_13_state_state <= _GEN_992;
                end
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_state_state <= 2'h0;
                end else begin
                  TBEMemory_13_state_state <= _GEN_992;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_13_state_state <= _GEN_992;
                end else if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_13_state_state <= _GEN_992;
                end
              end else begin
                TBEMemory_13_state_state <= _GEN_992;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEMemory_13_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_13_state_state <= _GEN_992;
                  end
                end else if (_T_133) begin
                  if (4'hd == idxUpdate_2[3:0]) begin
                    TBEMemory_13_state_state <= 2'h0;
                  end else begin
                    TBEMemory_13_state_state <= _GEN_992;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_13_state_state <= _GEN_992;
                  end else if (4'hd == idxUpdate_2[3:0]) begin
                    TBEMemory_13_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_13_state_state <= _GEN_992;
                  end
                end else begin
                  TBEMemory_13_state_state <= _GEN_992;
                end
              end else if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEMemory_13_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_13_state_state <= _GEN_992;
                end
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_state_state <= 2'h0;
                end else begin
                  TBEMemory_13_state_state <= _GEN_992;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_13_state_state <= _GEN_992;
                end else if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_13_state_state <= _GEN_992;
                end
              end else begin
                TBEMemory_13_state_state <= _GEN_992;
              end
            end else begin
              TBEMemory_13_state_state <= _GEN_1506;
            end
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEMemory_13_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_13_state_state <= _GEN_1506;
              end
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_state_state <= 2'h0;
              end else begin
                TBEMemory_13_state_state <= _GEN_1506;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_13_state_state <= _GEN_1506;
              end else if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_13_state_state <= _GEN_1506;
              end
            end else begin
              TBEMemory_13_state_state <= _GEN_1506;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEMemory_13_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_13_state_state <= _GEN_1506;
                end
              end else if (_T_155) begin
                if (4'hd == idxUpdate_3[3:0]) begin
                  TBEMemory_13_state_state <= 2'h0;
                end else begin
                  TBEMemory_13_state_state <= _GEN_1506;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_13_state_state <= _GEN_1506;
                end else if (4'hd == idxUpdate_3[3:0]) begin
                  TBEMemory_13_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_13_state_state <= _GEN_1506;
                end
              end else begin
                TBEMemory_13_state_state <= _GEN_1506;
              end
            end else if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEMemory_13_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_13_state_state <= _GEN_1506;
              end
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_state_state <= 2'h0;
              end else begin
                TBEMemory_13_state_state <= _GEN_1506;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_13_state_state <= _GEN_1506;
              end else if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_13_state_state <= _GEN_1506;
              end
            end else begin
              TBEMemory_13_state_state <= _GEN_1506;
            end
          end else begin
            TBEMemory_13_state_state <= _GEN_2020;
          end
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEMemory_13_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_13_state_state <= _GEN_2020;
            end
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_state_state <= 2'h0;
            end else begin
              TBEMemory_13_state_state <= _GEN_2020;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_13_state_state <= _GEN_2020;
            end else if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_13_state_state <= _GEN_2020;
            end
          end else begin
            TBEMemory_13_state_state <= _GEN_2020;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEMemory_13_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_13_state_state <= _GEN_2020;
              end
            end else if (_T_177) begin
              if (4'hd == idxUpdate_4[3:0]) begin
                TBEMemory_13_state_state <= 2'h0;
              end else begin
                TBEMemory_13_state_state <= _GEN_2020;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_13_state_state <= _GEN_2020;
              end else if (4'hd == idxUpdate_4[3:0]) begin
                TBEMemory_13_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_13_state_state <= _GEN_2020;
              end
            end else begin
              TBEMemory_13_state_state <= _GEN_2020;
            end
          end else if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEMemory_13_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_13_state_state <= _GEN_2020;
            end
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_state_state <= 2'h0;
            end else begin
              TBEMemory_13_state_state <= _GEN_2020;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_13_state_state <= _GEN_2020;
            end else if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_13_state_state <= _GEN_2020;
            end
          end else begin
            TBEMemory_13_state_state <= _GEN_2020;
          end
        end else begin
          TBEMemory_13_state_state <= _GEN_2534;
        end
      end else if (_T_221) begin
        if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEMemory_13_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_13_state_state <= _GEN_2534;
          end
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_state_state <= 2'h0;
          end else begin
            TBEMemory_13_state_state <= _GEN_2534;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_13_state_state <= _GEN_2534;
          end else if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_13_state_state <= _GEN_2534;
          end
        end else begin
          TBEMemory_13_state_state <= _GEN_2534;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEMemory_13_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_13_state_state <= _GEN_2534;
            end
          end else if (_T_199) begin
            if (4'hd == idxUpdate_5[3:0]) begin
              TBEMemory_13_state_state <= 2'h0;
            end else begin
              TBEMemory_13_state_state <= _GEN_2534;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_13_state_state <= _GEN_2534;
            end else if (4'hd == idxUpdate_5[3:0]) begin
              TBEMemory_13_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_13_state_state <= _GEN_2534;
            end
          end else begin
            TBEMemory_13_state_state <= _GEN_2534;
          end
        end else if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEMemory_13_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_13_state_state <= _GEN_2534;
          end
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_state_state <= 2'h0;
          end else begin
            TBEMemory_13_state_state <= _GEN_2534;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_13_state_state <= _GEN_2534;
          end else if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_13_state_state <= _GEN_2534;
          end
        end else begin
          TBEMemory_13_state_state <= _GEN_2534;
        end
      end else begin
        TBEMemory_13_state_state <= _GEN_3048;
      end
    end else if (_T_243) begin
      if (4'hd == idxUpdate_7[3:0]) begin
        TBEMemory_13_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'hd == idxAlloc[3:0]) begin
          TBEMemory_13_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_13_state_state <= _GEN_3048;
        end
      end else if (_T_221) begin
        if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_state_state <= 2'h0;
        end else begin
          TBEMemory_13_state_state <= _GEN_3048;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_13_state_state <= _GEN_3048;
        end else if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_13_state_state <= _GEN_3048;
        end
      end else begin
        TBEMemory_13_state_state <= _GEN_3048;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEMemory_13_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_13_state_state <= _GEN_3048;
          end
        end else if (_T_221) begin
          if (4'hd == idxUpdate_6[3:0]) begin
            TBEMemory_13_state_state <= 2'h0;
          end else begin
            TBEMemory_13_state_state <= _GEN_3048;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_13_state_state <= _GEN_3048;
          end else if (4'hd == idxUpdate_6[3:0]) begin
            TBEMemory_13_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_13_state_state <= _GEN_3048;
          end
        end else begin
          TBEMemory_13_state_state <= _GEN_3048;
        end
      end else if (4'hd == idxUpdate_7[3:0]) begin
        TBEMemory_13_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'hd == idxAlloc[3:0]) begin
          TBEMemory_13_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_13_state_state <= _GEN_3048;
        end
      end else if (_T_221) begin
        if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_state_state <= 2'h0;
        end else begin
          TBEMemory_13_state_state <= _GEN_3048;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_13_state_state <= _GEN_3048;
        end else if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_13_state_state <= _GEN_3048;
        end
      end else begin
        TBEMemory_13_state_state <= _GEN_3048;
      end
    end else begin
      TBEMemory_13_state_state <= _GEN_3562;
    end
    if (reset) begin
      TBEMemory_13_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'hd == idxAlloc[3:0]) begin
        TBEMemory_13_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'hd == idxAlloc[3:0]) begin
          TBEMemory_13_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEMemory_13_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEMemory_13_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEMemory_13_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEMemory_13_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEMemory_13_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEMemory_13_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEMemory_13_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hd == idxUpdate_0[3:0]) begin
                        TBEMemory_13_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEMemory_13_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEMemory_13_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hd == idxUpdate_0[3:0]) begin
                        TBEMemory_13_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'hd == idxAlloc[3:0]) begin
                        TBEMemory_13_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'hd == idxUpdate_0[3:0]) begin
                        TBEMemory_13_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'hd == idxUpdate_0[3:0]) begin
                          TBEMemory_13_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEMemory_13_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEMemory_13_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hd == idxUpdate_0[3:0]) begin
                        TBEMemory_13_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_13_way <= _GEN_462;
                end
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEMemory_13_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_13_way <= _GEN_462;
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_way <= 3'h2;
                  end else begin
                    TBEMemory_13_way <= _GEN_462;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_13_way <= _GEN_462;
                  end else if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_13_way <= _GEN_462;
                  end
                end else begin
                  TBEMemory_13_way <= _GEN_462;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEMemory_13_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_13_way <= _GEN_462;
                    end
                  end else if (_T_111) begin
                    if (4'hd == idxUpdate_1[3:0]) begin
                      TBEMemory_13_way <= 3'h2;
                    end else begin
                      TBEMemory_13_way <= _GEN_462;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_13_way <= _GEN_462;
                    end else if (4'hd == idxUpdate_1[3:0]) begin
                      TBEMemory_13_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_13_way <= _GEN_462;
                    end
                  end else begin
                    TBEMemory_13_way <= _GEN_462;
                  end
                end else if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEMemory_13_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_13_way <= _GEN_462;
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_way <= 3'h2;
                  end else begin
                    TBEMemory_13_way <= _GEN_462;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_13_way <= _GEN_462;
                  end else if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_13_way <= _GEN_462;
                  end
                end else begin
                  TBEMemory_13_way <= _GEN_462;
                end
              end else begin
                TBEMemory_13_way <= _GEN_976;
              end
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEMemory_13_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_13_way <= _GEN_976;
                end
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_way <= 3'h2;
                end else begin
                  TBEMemory_13_way <= _GEN_976;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_13_way <= _GEN_976;
                end else if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_13_way <= _GEN_976;
                end
              end else begin
                TBEMemory_13_way <= _GEN_976;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEMemory_13_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_13_way <= _GEN_976;
                  end
                end else if (_T_133) begin
                  if (4'hd == idxUpdate_2[3:0]) begin
                    TBEMemory_13_way <= 3'h2;
                  end else begin
                    TBEMemory_13_way <= _GEN_976;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_13_way <= _GEN_976;
                  end else if (4'hd == idxUpdate_2[3:0]) begin
                    TBEMemory_13_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_13_way <= _GEN_976;
                  end
                end else begin
                  TBEMemory_13_way <= _GEN_976;
                end
              end else if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEMemory_13_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_13_way <= _GEN_976;
                end
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_way <= 3'h2;
                end else begin
                  TBEMemory_13_way <= _GEN_976;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_13_way <= _GEN_976;
                end else if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_13_way <= _GEN_976;
                end
              end else begin
                TBEMemory_13_way <= _GEN_976;
              end
            end else begin
              TBEMemory_13_way <= _GEN_1490;
            end
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEMemory_13_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_13_way <= _GEN_1490;
              end
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_way <= 3'h2;
              end else begin
                TBEMemory_13_way <= _GEN_1490;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_13_way <= _GEN_1490;
              end else if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_13_way <= _GEN_1490;
              end
            end else begin
              TBEMemory_13_way <= _GEN_1490;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEMemory_13_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_13_way <= _GEN_1490;
                end
              end else if (_T_155) begin
                if (4'hd == idxUpdate_3[3:0]) begin
                  TBEMemory_13_way <= 3'h2;
                end else begin
                  TBEMemory_13_way <= _GEN_1490;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_13_way <= _GEN_1490;
                end else if (4'hd == idxUpdate_3[3:0]) begin
                  TBEMemory_13_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_13_way <= _GEN_1490;
                end
              end else begin
                TBEMemory_13_way <= _GEN_1490;
              end
            end else if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEMemory_13_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_13_way <= _GEN_1490;
              end
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_way <= 3'h2;
              end else begin
                TBEMemory_13_way <= _GEN_1490;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_13_way <= _GEN_1490;
              end else if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_13_way <= _GEN_1490;
              end
            end else begin
              TBEMemory_13_way <= _GEN_1490;
            end
          end else begin
            TBEMemory_13_way <= _GEN_2004;
          end
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEMemory_13_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_13_way <= _GEN_2004;
            end
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_way <= 3'h2;
            end else begin
              TBEMemory_13_way <= _GEN_2004;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_13_way <= _GEN_2004;
            end else if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_13_way <= _GEN_2004;
            end
          end else begin
            TBEMemory_13_way <= _GEN_2004;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEMemory_13_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_13_way <= _GEN_2004;
              end
            end else if (_T_177) begin
              if (4'hd == idxUpdate_4[3:0]) begin
                TBEMemory_13_way <= 3'h2;
              end else begin
                TBEMemory_13_way <= _GEN_2004;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_13_way <= _GEN_2004;
              end else if (4'hd == idxUpdate_4[3:0]) begin
                TBEMemory_13_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_13_way <= _GEN_2004;
              end
            end else begin
              TBEMemory_13_way <= _GEN_2004;
            end
          end else if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEMemory_13_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_13_way <= _GEN_2004;
            end
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_way <= 3'h2;
            end else begin
              TBEMemory_13_way <= _GEN_2004;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_13_way <= _GEN_2004;
            end else if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_13_way <= _GEN_2004;
            end
          end else begin
            TBEMemory_13_way <= _GEN_2004;
          end
        end else begin
          TBEMemory_13_way <= _GEN_2518;
        end
      end else if (_T_221) begin
        if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEMemory_13_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_13_way <= _GEN_2518;
          end
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_way <= 3'h2;
          end else begin
            TBEMemory_13_way <= _GEN_2518;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_13_way <= _GEN_2518;
          end else if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_13_way <= _GEN_2518;
          end
        end else begin
          TBEMemory_13_way <= _GEN_2518;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEMemory_13_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_13_way <= _GEN_2518;
            end
          end else if (_T_199) begin
            if (4'hd == idxUpdate_5[3:0]) begin
              TBEMemory_13_way <= 3'h2;
            end else begin
              TBEMemory_13_way <= _GEN_2518;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_13_way <= _GEN_2518;
            end else if (4'hd == idxUpdate_5[3:0]) begin
              TBEMemory_13_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_13_way <= _GEN_2518;
            end
          end else begin
            TBEMemory_13_way <= _GEN_2518;
          end
        end else if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEMemory_13_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_13_way <= _GEN_2518;
          end
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_way <= 3'h2;
          end else begin
            TBEMemory_13_way <= _GEN_2518;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_13_way <= _GEN_2518;
          end else if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_13_way <= _GEN_2518;
          end
        end else begin
          TBEMemory_13_way <= _GEN_2518;
        end
      end else begin
        TBEMemory_13_way <= _GEN_3032;
      end
    end else if (_T_243) begin
      if (4'hd == idxUpdate_7[3:0]) begin
        TBEMemory_13_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'hd == idxAlloc[3:0]) begin
          TBEMemory_13_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_13_way <= _GEN_3032;
        end
      end else if (_T_221) begin
        if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_way <= 3'h2;
        end else begin
          TBEMemory_13_way <= _GEN_3032;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_13_way <= _GEN_3032;
        end else if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_13_way <= _GEN_3032;
        end
      end else begin
        TBEMemory_13_way <= _GEN_3032;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEMemory_13_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_13_way <= _GEN_3032;
          end
        end else if (_T_221) begin
          if (4'hd == idxUpdate_6[3:0]) begin
            TBEMemory_13_way <= 3'h2;
          end else begin
            TBEMemory_13_way <= _GEN_3032;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_13_way <= _GEN_3032;
          end else if (4'hd == idxUpdate_6[3:0]) begin
            TBEMemory_13_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_13_way <= _GEN_3032;
          end
        end else begin
          TBEMemory_13_way <= _GEN_3032;
        end
      end else if (4'hd == idxUpdate_7[3:0]) begin
        TBEMemory_13_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'hd == idxAlloc[3:0]) begin
          TBEMemory_13_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_13_way <= _GEN_3032;
        end
      end else if (_T_221) begin
        if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_way <= 3'h2;
        end else begin
          TBEMemory_13_way <= _GEN_3032;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_13_way <= _GEN_3032;
        end else if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_13_way <= _GEN_3032;
        end
      end else begin
        TBEMemory_13_way <= _GEN_3032;
      end
    end else begin
      TBEMemory_13_way <= _GEN_3546;
    end
    if (reset) begin
      TBEMemory_13_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'hd == idxAlloc[3:0]) begin
        TBEMemory_13_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'hd == idxAlloc[3:0]) begin
          TBEMemory_13_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEMemory_13_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEMemory_13_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEMemory_13_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEMemory_13_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEMemory_13_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEMemory_13_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEMemory_13_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'hd == idxUpdate_0[3:0]) begin
                        TBEMemory_13_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEMemory_13_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEMemory_13_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'hd == idxUpdate_0[3:0]) begin
                        TBEMemory_13_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'hd == idxUpdate_1[3:0]) begin
                      TBEMemory_13_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'hd == idxAlloc[3:0]) begin
                        TBEMemory_13_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'hd == idxUpdate_0[3:0]) begin
                        TBEMemory_13_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'hd == idxUpdate_0[3:0]) begin
                          TBEMemory_13_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEMemory_13_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEMemory_13_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'hd == idxUpdate_0[3:0]) begin
                        TBEMemory_13_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_446;
                end
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEMemory_13_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_446;
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_446;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'hd == idxUpdate_1[3:0]) begin
                      TBEMemory_13_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_13_fields_0 <= _GEN_446;
                    end
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_446;
                  end
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_446;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'hd == idxUpdate_2[3:0]) begin
                    TBEMemory_13_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEMemory_13_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_13_fields_0 <= _GEN_446;
                    end
                  end else if (_T_111) begin
                    if (4'hd == idxUpdate_1[3:0]) begin
                      TBEMemory_13_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_13_fields_0 <= _GEN_446;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'hd == idxUpdate_1[3:0]) begin
                        TBEMemory_13_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_13_fields_0 <= _GEN_446;
                      end
                    end else begin
                      TBEMemory_13_fields_0 <= _GEN_446;
                    end
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_446;
                  end
                end else if (isAlloc_1) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEMemory_13_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_446;
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEMemory_13_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_446;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'hd == idxUpdate_1[3:0]) begin
                      TBEMemory_13_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_13_fields_0 <= _GEN_446;
                    end
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_446;
                  end
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_446;
                end
              end else begin
                TBEMemory_13_fields_0 <= _GEN_960;
              end
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEMemory_13_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_960;
                end
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_960;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'hd == idxUpdate_2[3:0]) begin
                    TBEMemory_13_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_960;
                  end
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_960;
                end
              end else begin
                TBEMemory_13_fields_0 <= _GEN_960;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'hd == idxUpdate_3[3:0]) begin
                  TBEMemory_13_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEMemory_13_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_960;
                  end
                end else if (_T_133) begin
                  if (4'hd == idxUpdate_2[3:0]) begin
                    TBEMemory_13_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_960;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'hd == idxUpdate_2[3:0]) begin
                      TBEMemory_13_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_13_fields_0 <= _GEN_960;
                    end
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_960;
                  end
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_960;
                end
              end else if (isAlloc_2) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEMemory_13_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_960;
                end
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEMemory_13_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_960;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'hd == idxUpdate_2[3:0]) begin
                    TBEMemory_13_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_960;
                  end
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_960;
                end
              end else begin
                TBEMemory_13_fields_0 <= _GEN_960;
              end
            end else begin
              TBEMemory_13_fields_0 <= _GEN_1474;
            end
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEMemory_13_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_13_fields_0 <= _GEN_1474;
              end
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_fields_0 <= 32'h0;
              end else begin
                TBEMemory_13_fields_0 <= _GEN_1474;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'hd == idxUpdate_3[3:0]) begin
                  TBEMemory_13_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_1474;
                end
              end else begin
                TBEMemory_13_fields_0 <= _GEN_1474;
              end
            end else begin
              TBEMemory_13_fields_0 <= _GEN_1474;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'hd == idxUpdate_4[3:0]) begin
                TBEMemory_13_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEMemory_13_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_1474;
                end
              end else if (_T_155) begin
                if (4'hd == idxUpdate_3[3:0]) begin
                  TBEMemory_13_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_1474;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'hd == idxUpdate_3[3:0]) begin
                    TBEMemory_13_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_13_fields_0 <= _GEN_1474;
                  end
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_1474;
                end
              end else begin
                TBEMemory_13_fields_0 <= _GEN_1474;
              end
            end else if (isAlloc_3) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEMemory_13_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_13_fields_0 <= _GEN_1474;
              end
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEMemory_13_fields_0 <= 32'h0;
              end else begin
                TBEMemory_13_fields_0 <= _GEN_1474;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'hd == idxUpdate_3[3:0]) begin
                  TBEMemory_13_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_1474;
                end
              end else begin
                TBEMemory_13_fields_0 <= _GEN_1474;
              end
            end else begin
              TBEMemory_13_fields_0 <= _GEN_1474;
            end
          end else begin
            TBEMemory_13_fields_0 <= _GEN_1988;
          end
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEMemory_13_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_13_fields_0 <= _GEN_1988;
            end
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_fields_0 <= 32'h0;
            end else begin
              TBEMemory_13_fields_0 <= _GEN_1988;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'hd == idxUpdate_4[3:0]) begin
                TBEMemory_13_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_13_fields_0 <= _GEN_1988;
              end
            end else begin
              TBEMemory_13_fields_0 <= _GEN_1988;
            end
          end else begin
            TBEMemory_13_fields_0 <= _GEN_1988;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'hd == idxUpdate_5[3:0]) begin
              TBEMemory_13_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEMemory_13_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_13_fields_0 <= _GEN_1988;
              end
            end else if (_T_177) begin
              if (4'hd == idxUpdate_4[3:0]) begin
                TBEMemory_13_fields_0 <= 32'h0;
              end else begin
                TBEMemory_13_fields_0 <= _GEN_1988;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'hd == idxUpdate_4[3:0]) begin
                  TBEMemory_13_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_13_fields_0 <= _GEN_1988;
                end
              end else begin
                TBEMemory_13_fields_0 <= _GEN_1988;
              end
            end else begin
              TBEMemory_13_fields_0 <= _GEN_1988;
            end
          end else if (isAlloc_4) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEMemory_13_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_13_fields_0 <= _GEN_1988;
            end
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEMemory_13_fields_0 <= 32'h0;
            end else begin
              TBEMemory_13_fields_0 <= _GEN_1988;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'hd == idxUpdate_4[3:0]) begin
                TBEMemory_13_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_13_fields_0 <= _GEN_1988;
              end
            end else begin
              TBEMemory_13_fields_0 <= _GEN_1988;
            end
          end else begin
            TBEMemory_13_fields_0 <= _GEN_1988;
          end
        end else begin
          TBEMemory_13_fields_0 <= _GEN_2502;
        end
      end else if (_T_221) begin
        if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEMemory_13_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_13_fields_0 <= _GEN_2502;
          end
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_fields_0 <= 32'h0;
          end else begin
            TBEMemory_13_fields_0 <= _GEN_2502;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'hd == idxUpdate_5[3:0]) begin
              TBEMemory_13_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_13_fields_0 <= _GEN_2502;
            end
          end else begin
            TBEMemory_13_fields_0 <= _GEN_2502;
          end
        end else begin
          TBEMemory_13_fields_0 <= _GEN_2502;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'hd == idxUpdate_6[3:0]) begin
            TBEMemory_13_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEMemory_13_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_13_fields_0 <= _GEN_2502;
            end
          end else if (_T_199) begin
            if (4'hd == idxUpdate_5[3:0]) begin
              TBEMemory_13_fields_0 <= 32'h0;
            end else begin
              TBEMemory_13_fields_0 <= _GEN_2502;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'hd == idxUpdate_5[3:0]) begin
                TBEMemory_13_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_13_fields_0 <= _GEN_2502;
              end
            end else begin
              TBEMemory_13_fields_0 <= _GEN_2502;
            end
          end else begin
            TBEMemory_13_fields_0 <= _GEN_2502;
          end
        end else if (isAlloc_5) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEMemory_13_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_13_fields_0 <= _GEN_2502;
          end
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEMemory_13_fields_0 <= 32'h0;
          end else begin
            TBEMemory_13_fields_0 <= _GEN_2502;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'hd == idxUpdate_5[3:0]) begin
              TBEMemory_13_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_13_fields_0 <= _GEN_2502;
            end
          end else begin
            TBEMemory_13_fields_0 <= _GEN_2502;
          end
        end else begin
          TBEMemory_13_fields_0 <= _GEN_2502;
        end
      end else begin
        TBEMemory_13_fields_0 <= _GEN_3016;
      end
    end else if (_T_243) begin
      if (4'hd == idxUpdate_7[3:0]) begin
        TBEMemory_13_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'hd == idxAlloc[3:0]) begin
          TBEMemory_13_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_13_fields_0 <= _GEN_3016;
        end
      end else if (_T_221) begin
        if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_fields_0 <= 32'h0;
        end else begin
          TBEMemory_13_fields_0 <= _GEN_3016;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'hd == idxUpdate_6[3:0]) begin
            TBEMemory_13_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_13_fields_0 <= _GEN_3016;
          end
        end else begin
          TBEMemory_13_fields_0 <= _GEN_3016;
        end
      end else begin
        TBEMemory_13_fields_0 <= _GEN_3016;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'hd == idxUpdate_7[3:0]) begin
          TBEMemory_13_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEMemory_13_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_13_fields_0 <= _GEN_3016;
          end
        end else if (_T_221) begin
          if (4'hd == idxUpdate_6[3:0]) begin
            TBEMemory_13_fields_0 <= 32'h0;
          end else begin
            TBEMemory_13_fields_0 <= _GEN_3016;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'hd == idxUpdate_6[3:0]) begin
              TBEMemory_13_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_13_fields_0 <= _GEN_3016;
            end
          end else begin
            TBEMemory_13_fields_0 <= _GEN_3016;
          end
        end else begin
          TBEMemory_13_fields_0 <= _GEN_3016;
        end
      end else if (isAlloc_6) begin
        if (4'hd == idxAlloc[3:0]) begin
          TBEMemory_13_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_13_fields_0 <= _GEN_3016;
        end
      end else if (_T_221) begin
        if (4'hd == idxUpdate_6[3:0]) begin
          TBEMemory_13_fields_0 <= 32'h0;
        end else begin
          TBEMemory_13_fields_0 <= _GEN_3016;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'hd == idxUpdate_6[3:0]) begin
            TBEMemory_13_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_13_fields_0 <= _GEN_3016;
          end
        end else begin
          TBEMemory_13_fields_0 <= _GEN_3016;
        end
      end else begin
        TBEMemory_13_fields_0 <= _GEN_3016;
      end
    end else begin
      TBEMemory_13_fields_0 <= _GEN_3530;
    end
    if (reset) begin
      TBEMemory_14_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'he == idxAlloc[3:0]) begin
        TBEMemory_14_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'he == idxAlloc[3:0]) begin
          TBEMemory_14_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEMemory_14_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEMemory_14_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEMemory_14_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEMemory_14_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEMemory_14_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEMemory_14_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEMemory_14_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'he == idxUpdate_0[3:0]) begin
                        TBEMemory_14_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEMemory_14_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEMemory_14_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'he == idxUpdate_0[3:0]) begin
                        TBEMemory_14_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'he == idxAlloc[3:0]) begin
                        TBEMemory_14_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'he == idxUpdate_0[3:0]) begin
                        TBEMemory_14_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'he == idxUpdate_0[3:0]) begin
                          TBEMemory_14_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEMemory_14_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEMemory_14_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'he == idxUpdate_0[3:0]) begin
                        TBEMemory_14_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_14_state_state <= _GEN_479;
                end
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEMemory_14_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_14_state_state <= _GEN_479;
                  end
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_state_state <= 2'h0;
                  end else begin
                    TBEMemory_14_state_state <= _GEN_479;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_14_state_state <= _GEN_479;
                  end else if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_14_state_state <= _GEN_479;
                  end
                end else begin
                  TBEMemory_14_state_state <= _GEN_479;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEMemory_14_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_14_state_state <= _GEN_479;
                    end
                  end else if (_T_111) begin
                    if (4'he == idxUpdate_1[3:0]) begin
                      TBEMemory_14_state_state <= 2'h0;
                    end else begin
                      TBEMemory_14_state_state <= _GEN_479;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_14_state_state <= _GEN_479;
                    end else if (4'he == idxUpdate_1[3:0]) begin
                      TBEMemory_14_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_14_state_state <= _GEN_479;
                    end
                  end else begin
                    TBEMemory_14_state_state <= _GEN_479;
                  end
                end else if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEMemory_14_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_14_state_state <= _GEN_479;
                  end
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_state_state <= 2'h0;
                  end else begin
                    TBEMemory_14_state_state <= _GEN_479;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_14_state_state <= _GEN_479;
                  end else if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_14_state_state <= _GEN_479;
                  end
                end else begin
                  TBEMemory_14_state_state <= _GEN_479;
                end
              end else begin
                TBEMemory_14_state_state <= _GEN_993;
              end
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEMemory_14_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_14_state_state <= _GEN_993;
                end
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_state_state <= 2'h0;
                end else begin
                  TBEMemory_14_state_state <= _GEN_993;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_14_state_state <= _GEN_993;
                end else if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_14_state_state <= _GEN_993;
                end
              end else begin
                TBEMemory_14_state_state <= _GEN_993;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEMemory_14_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_14_state_state <= _GEN_993;
                  end
                end else if (_T_133) begin
                  if (4'he == idxUpdate_2[3:0]) begin
                    TBEMemory_14_state_state <= 2'h0;
                  end else begin
                    TBEMemory_14_state_state <= _GEN_993;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_14_state_state <= _GEN_993;
                  end else if (4'he == idxUpdate_2[3:0]) begin
                    TBEMemory_14_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_14_state_state <= _GEN_993;
                  end
                end else begin
                  TBEMemory_14_state_state <= _GEN_993;
                end
              end else if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEMemory_14_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_14_state_state <= _GEN_993;
                end
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_state_state <= 2'h0;
                end else begin
                  TBEMemory_14_state_state <= _GEN_993;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_14_state_state <= _GEN_993;
                end else if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_14_state_state <= _GEN_993;
                end
              end else begin
                TBEMemory_14_state_state <= _GEN_993;
              end
            end else begin
              TBEMemory_14_state_state <= _GEN_1507;
            end
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEMemory_14_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_14_state_state <= _GEN_1507;
              end
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_state_state <= 2'h0;
              end else begin
                TBEMemory_14_state_state <= _GEN_1507;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_14_state_state <= _GEN_1507;
              end else if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_14_state_state <= _GEN_1507;
              end
            end else begin
              TBEMemory_14_state_state <= _GEN_1507;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEMemory_14_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_14_state_state <= _GEN_1507;
                end
              end else if (_T_155) begin
                if (4'he == idxUpdate_3[3:0]) begin
                  TBEMemory_14_state_state <= 2'h0;
                end else begin
                  TBEMemory_14_state_state <= _GEN_1507;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_14_state_state <= _GEN_1507;
                end else if (4'he == idxUpdate_3[3:0]) begin
                  TBEMemory_14_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_14_state_state <= _GEN_1507;
                end
              end else begin
                TBEMemory_14_state_state <= _GEN_1507;
              end
            end else if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEMemory_14_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_14_state_state <= _GEN_1507;
              end
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_state_state <= 2'h0;
              end else begin
                TBEMemory_14_state_state <= _GEN_1507;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_14_state_state <= _GEN_1507;
              end else if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_14_state_state <= _GEN_1507;
              end
            end else begin
              TBEMemory_14_state_state <= _GEN_1507;
            end
          end else begin
            TBEMemory_14_state_state <= _GEN_2021;
          end
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEMemory_14_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_14_state_state <= _GEN_2021;
            end
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_state_state <= 2'h0;
            end else begin
              TBEMemory_14_state_state <= _GEN_2021;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_14_state_state <= _GEN_2021;
            end else if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_14_state_state <= _GEN_2021;
            end
          end else begin
            TBEMemory_14_state_state <= _GEN_2021;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEMemory_14_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_14_state_state <= _GEN_2021;
              end
            end else if (_T_177) begin
              if (4'he == idxUpdate_4[3:0]) begin
                TBEMemory_14_state_state <= 2'h0;
              end else begin
                TBEMemory_14_state_state <= _GEN_2021;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_14_state_state <= _GEN_2021;
              end else if (4'he == idxUpdate_4[3:0]) begin
                TBEMemory_14_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_14_state_state <= _GEN_2021;
              end
            end else begin
              TBEMemory_14_state_state <= _GEN_2021;
            end
          end else if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEMemory_14_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_14_state_state <= _GEN_2021;
            end
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_state_state <= 2'h0;
            end else begin
              TBEMemory_14_state_state <= _GEN_2021;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_14_state_state <= _GEN_2021;
            end else if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_14_state_state <= _GEN_2021;
            end
          end else begin
            TBEMemory_14_state_state <= _GEN_2021;
          end
        end else begin
          TBEMemory_14_state_state <= _GEN_2535;
        end
      end else if (_T_221) begin
        if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEMemory_14_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_14_state_state <= _GEN_2535;
          end
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_state_state <= 2'h0;
          end else begin
            TBEMemory_14_state_state <= _GEN_2535;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_14_state_state <= _GEN_2535;
          end else if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_14_state_state <= _GEN_2535;
          end
        end else begin
          TBEMemory_14_state_state <= _GEN_2535;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEMemory_14_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_14_state_state <= _GEN_2535;
            end
          end else if (_T_199) begin
            if (4'he == idxUpdate_5[3:0]) begin
              TBEMemory_14_state_state <= 2'h0;
            end else begin
              TBEMemory_14_state_state <= _GEN_2535;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_14_state_state <= _GEN_2535;
            end else if (4'he == idxUpdate_5[3:0]) begin
              TBEMemory_14_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_14_state_state <= _GEN_2535;
            end
          end else begin
            TBEMemory_14_state_state <= _GEN_2535;
          end
        end else if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEMemory_14_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_14_state_state <= _GEN_2535;
          end
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_state_state <= 2'h0;
          end else begin
            TBEMemory_14_state_state <= _GEN_2535;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_14_state_state <= _GEN_2535;
          end else if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_14_state_state <= _GEN_2535;
          end
        end else begin
          TBEMemory_14_state_state <= _GEN_2535;
        end
      end else begin
        TBEMemory_14_state_state <= _GEN_3049;
      end
    end else if (_T_243) begin
      if (4'he == idxUpdate_7[3:0]) begin
        TBEMemory_14_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'he == idxAlloc[3:0]) begin
          TBEMemory_14_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_14_state_state <= _GEN_3049;
        end
      end else if (_T_221) begin
        if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_state_state <= 2'h0;
        end else begin
          TBEMemory_14_state_state <= _GEN_3049;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_14_state_state <= _GEN_3049;
        end else if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_14_state_state <= _GEN_3049;
        end
      end else begin
        TBEMemory_14_state_state <= _GEN_3049;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEMemory_14_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_14_state_state <= _GEN_3049;
          end
        end else if (_T_221) begin
          if (4'he == idxUpdate_6[3:0]) begin
            TBEMemory_14_state_state <= 2'h0;
          end else begin
            TBEMemory_14_state_state <= _GEN_3049;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_14_state_state <= _GEN_3049;
          end else if (4'he == idxUpdate_6[3:0]) begin
            TBEMemory_14_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_14_state_state <= _GEN_3049;
          end
        end else begin
          TBEMemory_14_state_state <= _GEN_3049;
        end
      end else if (4'he == idxUpdate_7[3:0]) begin
        TBEMemory_14_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'he == idxAlloc[3:0]) begin
          TBEMemory_14_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_14_state_state <= _GEN_3049;
        end
      end else if (_T_221) begin
        if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_state_state <= 2'h0;
        end else begin
          TBEMemory_14_state_state <= _GEN_3049;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_14_state_state <= _GEN_3049;
        end else if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_14_state_state <= _GEN_3049;
        end
      end else begin
        TBEMemory_14_state_state <= _GEN_3049;
      end
    end else begin
      TBEMemory_14_state_state <= _GEN_3563;
    end
    if (reset) begin
      TBEMemory_14_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'he == idxAlloc[3:0]) begin
        TBEMemory_14_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'he == idxAlloc[3:0]) begin
          TBEMemory_14_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEMemory_14_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEMemory_14_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEMemory_14_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEMemory_14_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEMemory_14_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEMemory_14_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEMemory_14_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'he == idxUpdate_0[3:0]) begin
                        TBEMemory_14_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEMemory_14_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEMemory_14_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'he == idxUpdate_0[3:0]) begin
                        TBEMemory_14_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'he == idxAlloc[3:0]) begin
                        TBEMemory_14_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'he == idxUpdate_0[3:0]) begin
                        TBEMemory_14_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'he == idxUpdate_0[3:0]) begin
                          TBEMemory_14_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEMemory_14_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEMemory_14_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'he == idxUpdate_0[3:0]) begin
                        TBEMemory_14_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_14_way <= _GEN_463;
                end
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEMemory_14_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_14_way <= _GEN_463;
                  end
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_way <= 3'h2;
                  end else begin
                    TBEMemory_14_way <= _GEN_463;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_14_way <= _GEN_463;
                  end else if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_14_way <= _GEN_463;
                  end
                end else begin
                  TBEMemory_14_way <= _GEN_463;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEMemory_14_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_14_way <= _GEN_463;
                    end
                  end else if (_T_111) begin
                    if (4'he == idxUpdate_1[3:0]) begin
                      TBEMemory_14_way <= 3'h2;
                    end else begin
                      TBEMemory_14_way <= _GEN_463;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_14_way <= _GEN_463;
                    end else if (4'he == idxUpdate_1[3:0]) begin
                      TBEMemory_14_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_14_way <= _GEN_463;
                    end
                  end else begin
                    TBEMemory_14_way <= _GEN_463;
                  end
                end else if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEMemory_14_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_14_way <= _GEN_463;
                  end
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_way <= 3'h2;
                  end else begin
                    TBEMemory_14_way <= _GEN_463;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_14_way <= _GEN_463;
                  end else if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_14_way <= _GEN_463;
                  end
                end else begin
                  TBEMemory_14_way <= _GEN_463;
                end
              end else begin
                TBEMemory_14_way <= _GEN_977;
              end
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEMemory_14_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_14_way <= _GEN_977;
                end
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_way <= 3'h2;
                end else begin
                  TBEMemory_14_way <= _GEN_977;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_14_way <= _GEN_977;
                end else if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_14_way <= _GEN_977;
                end
              end else begin
                TBEMemory_14_way <= _GEN_977;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEMemory_14_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_14_way <= _GEN_977;
                  end
                end else if (_T_133) begin
                  if (4'he == idxUpdate_2[3:0]) begin
                    TBEMemory_14_way <= 3'h2;
                  end else begin
                    TBEMemory_14_way <= _GEN_977;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_14_way <= _GEN_977;
                  end else if (4'he == idxUpdate_2[3:0]) begin
                    TBEMemory_14_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_14_way <= _GEN_977;
                  end
                end else begin
                  TBEMemory_14_way <= _GEN_977;
                end
              end else if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEMemory_14_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_14_way <= _GEN_977;
                end
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_way <= 3'h2;
                end else begin
                  TBEMemory_14_way <= _GEN_977;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_14_way <= _GEN_977;
                end else if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_14_way <= _GEN_977;
                end
              end else begin
                TBEMemory_14_way <= _GEN_977;
              end
            end else begin
              TBEMemory_14_way <= _GEN_1491;
            end
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEMemory_14_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_14_way <= _GEN_1491;
              end
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_way <= 3'h2;
              end else begin
                TBEMemory_14_way <= _GEN_1491;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_14_way <= _GEN_1491;
              end else if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_14_way <= _GEN_1491;
              end
            end else begin
              TBEMemory_14_way <= _GEN_1491;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEMemory_14_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_14_way <= _GEN_1491;
                end
              end else if (_T_155) begin
                if (4'he == idxUpdate_3[3:0]) begin
                  TBEMemory_14_way <= 3'h2;
                end else begin
                  TBEMemory_14_way <= _GEN_1491;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_14_way <= _GEN_1491;
                end else if (4'he == idxUpdate_3[3:0]) begin
                  TBEMemory_14_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_14_way <= _GEN_1491;
                end
              end else begin
                TBEMemory_14_way <= _GEN_1491;
              end
            end else if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEMemory_14_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_14_way <= _GEN_1491;
              end
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_way <= 3'h2;
              end else begin
                TBEMemory_14_way <= _GEN_1491;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_14_way <= _GEN_1491;
              end else if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_14_way <= _GEN_1491;
              end
            end else begin
              TBEMemory_14_way <= _GEN_1491;
            end
          end else begin
            TBEMemory_14_way <= _GEN_2005;
          end
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEMemory_14_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_14_way <= _GEN_2005;
            end
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_way <= 3'h2;
            end else begin
              TBEMemory_14_way <= _GEN_2005;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_14_way <= _GEN_2005;
            end else if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_14_way <= _GEN_2005;
            end
          end else begin
            TBEMemory_14_way <= _GEN_2005;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEMemory_14_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_14_way <= _GEN_2005;
              end
            end else if (_T_177) begin
              if (4'he == idxUpdate_4[3:0]) begin
                TBEMemory_14_way <= 3'h2;
              end else begin
                TBEMemory_14_way <= _GEN_2005;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_14_way <= _GEN_2005;
              end else if (4'he == idxUpdate_4[3:0]) begin
                TBEMemory_14_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_14_way <= _GEN_2005;
              end
            end else begin
              TBEMemory_14_way <= _GEN_2005;
            end
          end else if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEMemory_14_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_14_way <= _GEN_2005;
            end
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_way <= 3'h2;
            end else begin
              TBEMemory_14_way <= _GEN_2005;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_14_way <= _GEN_2005;
            end else if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_14_way <= _GEN_2005;
            end
          end else begin
            TBEMemory_14_way <= _GEN_2005;
          end
        end else begin
          TBEMemory_14_way <= _GEN_2519;
        end
      end else if (_T_221) begin
        if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEMemory_14_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_14_way <= _GEN_2519;
          end
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_way <= 3'h2;
          end else begin
            TBEMemory_14_way <= _GEN_2519;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_14_way <= _GEN_2519;
          end else if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_14_way <= _GEN_2519;
          end
        end else begin
          TBEMemory_14_way <= _GEN_2519;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEMemory_14_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_14_way <= _GEN_2519;
            end
          end else if (_T_199) begin
            if (4'he == idxUpdate_5[3:0]) begin
              TBEMemory_14_way <= 3'h2;
            end else begin
              TBEMemory_14_way <= _GEN_2519;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_14_way <= _GEN_2519;
            end else if (4'he == idxUpdate_5[3:0]) begin
              TBEMemory_14_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_14_way <= _GEN_2519;
            end
          end else begin
            TBEMemory_14_way <= _GEN_2519;
          end
        end else if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEMemory_14_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_14_way <= _GEN_2519;
          end
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_way <= 3'h2;
          end else begin
            TBEMemory_14_way <= _GEN_2519;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_14_way <= _GEN_2519;
          end else if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_14_way <= _GEN_2519;
          end
        end else begin
          TBEMemory_14_way <= _GEN_2519;
        end
      end else begin
        TBEMemory_14_way <= _GEN_3033;
      end
    end else if (_T_243) begin
      if (4'he == idxUpdate_7[3:0]) begin
        TBEMemory_14_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'he == idxAlloc[3:0]) begin
          TBEMemory_14_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_14_way <= _GEN_3033;
        end
      end else if (_T_221) begin
        if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_way <= 3'h2;
        end else begin
          TBEMemory_14_way <= _GEN_3033;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_14_way <= _GEN_3033;
        end else if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_14_way <= _GEN_3033;
        end
      end else begin
        TBEMemory_14_way <= _GEN_3033;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEMemory_14_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_14_way <= _GEN_3033;
          end
        end else if (_T_221) begin
          if (4'he == idxUpdate_6[3:0]) begin
            TBEMemory_14_way <= 3'h2;
          end else begin
            TBEMemory_14_way <= _GEN_3033;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_14_way <= _GEN_3033;
          end else if (4'he == idxUpdate_6[3:0]) begin
            TBEMemory_14_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_14_way <= _GEN_3033;
          end
        end else begin
          TBEMemory_14_way <= _GEN_3033;
        end
      end else if (4'he == idxUpdate_7[3:0]) begin
        TBEMemory_14_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'he == idxAlloc[3:0]) begin
          TBEMemory_14_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_14_way <= _GEN_3033;
        end
      end else if (_T_221) begin
        if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_way <= 3'h2;
        end else begin
          TBEMemory_14_way <= _GEN_3033;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_14_way <= _GEN_3033;
        end else if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_14_way <= _GEN_3033;
        end
      end else begin
        TBEMemory_14_way <= _GEN_3033;
      end
    end else begin
      TBEMemory_14_way <= _GEN_3547;
    end
    if (reset) begin
      TBEMemory_14_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'he == idxAlloc[3:0]) begin
        TBEMemory_14_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'he == idxAlloc[3:0]) begin
          TBEMemory_14_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEMemory_14_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEMemory_14_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEMemory_14_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEMemory_14_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEMemory_14_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEMemory_14_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEMemory_14_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'he == idxUpdate_0[3:0]) begin
                        TBEMemory_14_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEMemory_14_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEMemory_14_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'he == idxUpdate_0[3:0]) begin
                        TBEMemory_14_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'he == idxUpdate_1[3:0]) begin
                      TBEMemory_14_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'he == idxAlloc[3:0]) begin
                        TBEMemory_14_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'he == idxUpdate_0[3:0]) begin
                        TBEMemory_14_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'he == idxUpdate_0[3:0]) begin
                          TBEMemory_14_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEMemory_14_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEMemory_14_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'he == idxUpdate_0[3:0]) begin
                        TBEMemory_14_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_447;
                end
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEMemory_14_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_447;
                  end
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_447;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'he == idxUpdate_1[3:0]) begin
                      TBEMemory_14_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_14_fields_0 <= _GEN_447;
                    end
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_447;
                  end
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_447;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'he == idxUpdate_2[3:0]) begin
                    TBEMemory_14_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEMemory_14_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_14_fields_0 <= _GEN_447;
                    end
                  end else if (_T_111) begin
                    if (4'he == idxUpdate_1[3:0]) begin
                      TBEMemory_14_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_14_fields_0 <= _GEN_447;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'he == idxUpdate_1[3:0]) begin
                        TBEMemory_14_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_14_fields_0 <= _GEN_447;
                      end
                    end else begin
                      TBEMemory_14_fields_0 <= _GEN_447;
                    end
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_447;
                  end
                end else if (isAlloc_1) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEMemory_14_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_447;
                  end
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEMemory_14_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_447;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'he == idxUpdate_1[3:0]) begin
                      TBEMemory_14_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_14_fields_0 <= _GEN_447;
                    end
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_447;
                  end
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_447;
                end
              end else begin
                TBEMemory_14_fields_0 <= _GEN_961;
              end
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEMemory_14_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_961;
                end
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_961;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'he == idxUpdate_2[3:0]) begin
                    TBEMemory_14_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_961;
                  end
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_961;
                end
              end else begin
                TBEMemory_14_fields_0 <= _GEN_961;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'he == idxUpdate_3[3:0]) begin
                  TBEMemory_14_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEMemory_14_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_961;
                  end
                end else if (_T_133) begin
                  if (4'he == idxUpdate_2[3:0]) begin
                    TBEMemory_14_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_961;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'he == idxUpdate_2[3:0]) begin
                      TBEMemory_14_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_14_fields_0 <= _GEN_961;
                    end
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_961;
                  end
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_961;
                end
              end else if (isAlloc_2) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEMemory_14_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_961;
                end
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEMemory_14_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_961;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'he == idxUpdate_2[3:0]) begin
                    TBEMemory_14_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_961;
                  end
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_961;
                end
              end else begin
                TBEMemory_14_fields_0 <= _GEN_961;
              end
            end else begin
              TBEMemory_14_fields_0 <= _GEN_1475;
            end
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEMemory_14_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_14_fields_0 <= _GEN_1475;
              end
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_fields_0 <= 32'h0;
              end else begin
                TBEMemory_14_fields_0 <= _GEN_1475;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'he == idxUpdate_3[3:0]) begin
                  TBEMemory_14_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_1475;
                end
              end else begin
                TBEMemory_14_fields_0 <= _GEN_1475;
              end
            end else begin
              TBEMemory_14_fields_0 <= _GEN_1475;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'he == idxUpdate_4[3:0]) begin
                TBEMemory_14_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEMemory_14_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_1475;
                end
              end else if (_T_155) begin
                if (4'he == idxUpdate_3[3:0]) begin
                  TBEMemory_14_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_1475;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'he == idxUpdate_3[3:0]) begin
                    TBEMemory_14_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_14_fields_0 <= _GEN_1475;
                  end
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_1475;
                end
              end else begin
                TBEMemory_14_fields_0 <= _GEN_1475;
              end
            end else if (isAlloc_3) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEMemory_14_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_14_fields_0 <= _GEN_1475;
              end
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEMemory_14_fields_0 <= 32'h0;
              end else begin
                TBEMemory_14_fields_0 <= _GEN_1475;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'he == idxUpdate_3[3:0]) begin
                  TBEMemory_14_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_1475;
                end
              end else begin
                TBEMemory_14_fields_0 <= _GEN_1475;
              end
            end else begin
              TBEMemory_14_fields_0 <= _GEN_1475;
            end
          end else begin
            TBEMemory_14_fields_0 <= _GEN_1989;
          end
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEMemory_14_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_14_fields_0 <= _GEN_1989;
            end
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_fields_0 <= 32'h0;
            end else begin
              TBEMemory_14_fields_0 <= _GEN_1989;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'he == idxUpdate_4[3:0]) begin
                TBEMemory_14_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_14_fields_0 <= _GEN_1989;
              end
            end else begin
              TBEMemory_14_fields_0 <= _GEN_1989;
            end
          end else begin
            TBEMemory_14_fields_0 <= _GEN_1989;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'he == idxUpdate_5[3:0]) begin
              TBEMemory_14_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEMemory_14_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_14_fields_0 <= _GEN_1989;
              end
            end else if (_T_177) begin
              if (4'he == idxUpdate_4[3:0]) begin
                TBEMemory_14_fields_0 <= 32'h0;
              end else begin
                TBEMemory_14_fields_0 <= _GEN_1989;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'he == idxUpdate_4[3:0]) begin
                  TBEMemory_14_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_14_fields_0 <= _GEN_1989;
                end
              end else begin
                TBEMemory_14_fields_0 <= _GEN_1989;
              end
            end else begin
              TBEMemory_14_fields_0 <= _GEN_1989;
            end
          end else if (isAlloc_4) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEMemory_14_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_14_fields_0 <= _GEN_1989;
            end
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEMemory_14_fields_0 <= 32'h0;
            end else begin
              TBEMemory_14_fields_0 <= _GEN_1989;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'he == idxUpdate_4[3:0]) begin
                TBEMemory_14_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_14_fields_0 <= _GEN_1989;
              end
            end else begin
              TBEMemory_14_fields_0 <= _GEN_1989;
            end
          end else begin
            TBEMemory_14_fields_0 <= _GEN_1989;
          end
        end else begin
          TBEMemory_14_fields_0 <= _GEN_2503;
        end
      end else if (_T_221) begin
        if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEMemory_14_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_14_fields_0 <= _GEN_2503;
          end
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_fields_0 <= 32'h0;
          end else begin
            TBEMemory_14_fields_0 <= _GEN_2503;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'he == idxUpdate_5[3:0]) begin
              TBEMemory_14_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_14_fields_0 <= _GEN_2503;
            end
          end else begin
            TBEMemory_14_fields_0 <= _GEN_2503;
          end
        end else begin
          TBEMemory_14_fields_0 <= _GEN_2503;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'he == idxUpdate_6[3:0]) begin
            TBEMemory_14_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEMemory_14_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_14_fields_0 <= _GEN_2503;
            end
          end else if (_T_199) begin
            if (4'he == idxUpdate_5[3:0]) begin
              TBEMemory_14_fields_0 <= 32'h0;
            end else begin
              TBEMemory_14_fields_0 <= _GEN_2503;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'he == idxUpdate_5[3:0]) begin
                TBEMemory_14_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_14_fields_0 <= _GEN_2503;
              end
            end else begin
              TBEMemory_14_fields_0 <= _GEN_2503;
            end
          end else begin
            TBEMemory_14_fields_0 <= _GEN_2503;
          end
        end else if (isAlloc_5) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEMemory_14_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_14_fields_0 <= _GEN_2503;
          end
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEMemory_14_fields_0 <= 32'h0;
          end else begin
            TBEMemory_14_fields_0 <= _GEN_2503;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'he == idxUpdate_5[3:0]) begin
              TBEMemory_14_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_14_fields_0 <= _GEN_2503;
            end
          end else begin
            TBEMemory_14_fields_0 <= _GEN_2503;
          end
        end else begin
          TBEMemory_14_fields_0 <= _GEN_2503;
        end
      end else begin
        TBEMemory_14_fields_0 <= _GEN_3017;
      end
    end else if (_T_243) begin
      if (4'he == idxUpdate_7[3:0]) begin
        TBEMemory_14_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'he == idxAlloc[3:0]) begin
          TBEMemory_14_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_14_fields_0 <= _GEN_3017;
        end
      end else if (_T_221) begin
        if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_fields_0 <= 32'h0;
        end else begin
          TBEMemory_14_fields_0 <= _GEN_3017;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'he == idxUpdate_6[3:0]) begin
            TBEMemory_14_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_14_fields_0 <= _GEN_3017;
          end
        end else begin
          TBEMemory_14_fields_0 <= _GEN_3017;
        end
      end else begin
        TBEMemory_14_fields_0 <= _GEN_3017;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'he == idxUpdate_7[3:0]) begin
          TBEMemory_14_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEMemory_14_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_14_fields_0 <= _GEN_3017;
          end
        end else if (_T_221) begin
          if (4'he == idxUpdate_6[3:0]) begin
            TBEMemory_14_fields_0 <= 32'h0;
          end else begin
            TBEMemory_14_fields_0 <= _GEN_3017;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'he == idxUpdate_6[3:0]) begin
              TBEMemory_14_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_14_fields_0 <= _GEN_3017;
            end
          end else begin
            TBEMemory_14_fields_0 <= _GEN_3017;
          end
        end else begin
          TBEMemory_14_fields_0 <= _GEN_3017;
        end
      end else if (isAlloc_6) begin
        if (4'he == idxAlloc[3:0]) begin
          TBEMemory_14_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_14_fields_0 <= _GEN_3017;
        end
      end else if (_T_221) begin
        if (4'he == idxUpdate_6[3:0]) begin
          TBEMemory_14_fields_0 <= 32'h0;
        end else begin
          TBEMemory_14_fields_0 <= _GEN_3017;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'he == idxUpdate_6[3:0]) begin
            TBEMemory_14_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_14_fields_0 <= _GEN_3017;
          end
        end else begin
          TBEMemory_14_fields_0 <= _GEN_3017;
        end
      end else begin
        TBEMemory_14_fields_0 <= _GEN_3017;
      end
    end else begin
      TBEMemory_14_fields_0 <= _GEN_3531;
    end
    if (reset) begin
      TBEMemory_15_state_state <= 2'h0;
    end else if (isAlloc_7) begin
      if (4'hf == idxAlloc[3:0]) begin
        TBEMemory_15_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'hf == idxAlloc[3:0]) begin
          TBEMemory_15_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEMemory_15_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEMemory_15_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEMemory_15_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEMemory_15_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEMemory_15_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEMemory_15_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEMemory_15_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hf == idxUpdate_0[3:0]) begin
                        TBEMemory_15_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_state_state <= 2'h0;
                  end else if (isAlloc_0) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEMemory_15_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEMemory_15_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hf == idxUpdate_0[3:0]) begin
                        TBEMemory_15_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'hf == idxAlloc[3:0]) begin
                        TBEMemory_15_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end else if (_T_89) begin
                      if (4'hf == idxUpdate_0[3:0]) begin
                        TBEMemory_15_state_state <= 2'h0;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'hf == idxUpdate_0[3:0]) begin
                          TBEMemory_15_state_state <= io_write_0_bits_inputTBE_state_state;
                        end
                      end
                    end
                  end else if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else if (isAlloc_0) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEMemory_15_state_state <= io_write_0_bits_inputTBE_state_state;
                    end
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEMemory_15_state_state <= 2'h0;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hf == idxUpdate_0[3:0]) begin
                        TBEMemory_15_state_state <= io_write_0_bits_inputTBE_state_state;
                      end
                    end
                  end
                end else begin
                  TBEMemory_15_state_state <= _GEN_480;
                end
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_state_state <= 2'h0;
                end else if (isAlloc_1) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEMemory_15_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_15_state_state <= _GEN_480;
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_state_state <= 2'h0;
                  end else begin
                    TBEMemory_15_state_state <= _GEN_480;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_15_state_state <= _GEN_480;
                  end else if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_15_state_state <= _GEN_480;
                  end
                end else begin
                  TBEMemory_15_state_state <= _GEN_480;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEMemory_15_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_15_state_state <= _GEN_480;
                    end
                  end else if (_T_111) begin
                    if (4'hf == idxUpdate_1[3:0]) begin
                      TBEMemory_15_state_state <= 2'h0;
                    end else begin
                      TBEMemory_15_state_state <= _GEN_480;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_15_state_state <= _GEN_480;
                    end else if (4'hf == idxUpdate_1[3:0]) begin
                      TBEMemory_15_state_state <= io_write_1_bits_inputTBE_state_state;
                    end else begin
                      TBEMemory_15_state_state <= _GEN_480;
                    end
                  end else begin
                    TBEMemory_15_state_state <= _GEN_480;
                  end
                end else if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_state_state <= io_write_2_bits_inputTBE_state_state;
                end else if (isAlloc_1) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEMemory_15_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_15_state_state <= _GEN_480;
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_state_state <= 2'h0;
                  end else begin
                    TBEMemory_15_state_state <= _GEN_480;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_15_state_state <= _GEN_480;
                  end else if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_state_state <= io_write_1_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_15_state_state <= _GEN_480;
                  end
                end else begin
                  TBEMemory_15_state_state <= _GEN_480;
                end
              end else begin
                TBEMemory_15_state_state <= _GEN_994;
              end
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_state_state <= 2'h0;
              end else if (isAlloc_2) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEMemory_15_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_15_state_state <= _GEN_994;
                end
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_state_state <= 2'h0;
                end else begin
                  TBEMemory_15_state_state <= _GEN_994;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_15_state_state <= _GEN_994;
                end else if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_15_state_state <= _GEN_994;
                end
              end else begin
                TBEMemory_15_state_state <= _GEN_994;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEMemory_15_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_15_state_state <= _GEN_994;
                  end
                end else if (_T_133) begin
                  if (4'hf == idxUpdate_2[3:0]) begin
                    TBEMemory_15_state_state <= 2'h0;
                  end else begin
                    TBEMemory_15_state_state <= _GEN_994;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_15_state_state <= _GEN_994;
                  end else if (4'hf == idxUpdate_2[3:0]) begin
                    TBEMemory_15_state_state <= io_write_2_bits_inputTBE_state_state;
                  end else begin
                    TBEMemory_15_state_state <= _GEN_994;
                  end
                end else begin
                  TBEMemory_15_state_state <= _GEN_994;
                end
              end else if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_state_state <= io_write_3_bits_inputTBE_state_state;
              end else if (isAlloc_2) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEMemory_15_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_15_state_state <= _GEN_994;
                end
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_state_state <= 2'h0;
                end else begin
                  TBEMemory_15_state_state <= _GEN_994;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_15_state_state <= _GEN_994;
                end else if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_state_state <= io_write_2_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_15_state_state <= _GEN_994;
                end
              end else begin
                TBEMemory_15_state_state <= _GEN_994;
              end
            end else begin
              TBEMemory_15_state_state <= _GEN_1508;
            end
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_state_state <= 2'h0;
            end else if (isAlloc_3) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEMemory_15_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_15_state_state <= _GEN_1508;
              end
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_state_state <= 2'h0;
              end else begin
                TBEMemory_15_state_state <= _GEN_1508;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_15_state_state <= _GEN_1508;
              end else if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_15_state_state <= _GEN_1508;
              end
            end else begin
              TBEMemory_15_state_state <= _GEN_1508;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEMemory_15_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_15_state_state <= _GEN_1508;
                end
              end else if (_T_155) begin
                if (4'hf == idxUpdate_3[3:0]) begin
                  TBEMemory_15_state_state <= 2'h0;
                end else begin
                  TBEMemory_15_state_state <= _GEN_1508;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_15_state_state <= _GEN_1508;
                end else if (4'hf == idxUpdate_3[3:0]) begin
                  TBEMemory_15_state_state <= io_write_3_bits_inputTBE_state_state;
                end else begin
                  TBEMemory_15_state_state <= _GEN_1508;
                end
              end else begin
                TBEMemory_15_state_state <= _GEN_1508;
              end
            end else if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_state_state <= io_write_4_bits_inputTBE_state_state;
            end else if (isAlloc_3) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEMemory_15_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_15_state_state <= _GEN_1508;
              end
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_state_state <= 2'h0;
              end else begin
                TBEMemory_15_state_state <= _GEN_1508;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_15_state_state <= _GEN_1508;
              end else if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_state_state <= io_write_3_bits_inputTBE_state_state;
              end else begin
                TBEMemory_15_state_state <= _GEN_1508;
              end
            end else begin
              TBEMemory_15_state_state <= _GEN_1508;
            end
          end else begin
            TBEMemory_15_state_state <= _GEN_2022;
          end
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_state_state <= 2'h0;
          end else if (isAlloc_4) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEMemory_15_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_15_state_state <= _GEN_2022;
            end
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_state_state <= 2'h0;
            end else begin
              TBEMemory_15_state_state <= _GEN_2022;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_15_state_state <= _GEN_2022;
            end else if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_15_state_state <= _GEN_2022;
            end
          end else begin
            TBEMemory_15_state_state <= _GEN_2022;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEMemory_15_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_15_state_state <= _GEN_2022;
              end
            end else if (_T_177) begin
              if (4'hf == idxUpdate_4[3:0]) begin
                TBEMemory_15_state_state <= 2'h0;
              end else begin
                TBEMemory_15_state_state <= _GEN_2022;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_15_state_state <= _GEN_2022;
              end else if (4'hf == idxUpdate_4[3:0]) begin
                TBEMemory_15_state_state <= io_write_4_bits_inputTBE_state_state;
              end else begin
                TBEMemory_15_state_state <= _GEN_2022;
              end
            end else begin
              TBEMemory_15_state_state <= _GEN_2022;
            end
          end else if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_state_state <= io_write_5_bits_inputTBE_state_state;
          end else if (isAlloc_4) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEMemory_15_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_15_state_state <= _GEN_2022;
            end
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_state_state <= 2'h0;
            end else begin
              TBEMemory_15_state_state <= _GEN_2022;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_15_state_state <= _GEN_2022;
            end else if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_state_state <= io_write_4_bits_inputTBE_state_state;
            end else begin
              TBEMemory_15_state_state <= _GEN_2022;
            end
          end else begin
            TBEMemory_15_state_state <= _GEN_2022;
          end
        end else begin
          TBEMemory_15_state_state <= _GEN_2536;
        end
      end else if (_T_221) begin
        if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_state_state <= 2'h0;
        end else if (isAlloc_5) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEMemory_15_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_15_state_state <= _GEN_2536;
          end
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_state_state <= 2'h0;
          end else begin
            TBEMemory_15_state_state <= _GEN_2536;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_15_state_state <= _GEN_2536;
          end else if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_15_state_state <= _GEN_2536;
          end
        end else begin
          TBEMemory_15_state_state <= _GEN_2536;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEMemory_15_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_15_state_state <= _GEN_2536;
            end
          end else if (_T_199) begin
            if (4'hf == idxUpdate_5[3:0]) begin
              TBEMemory_15_state_state <= 2'h0;
            end else begin
              TBEMemory_15_state_state <= _GEN_2536;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_15_state_state <= _GEN_2536;
            end else if (4'hf == idxUpdate_5[3:0]) begin
              TBEMemory_15_state_state <= io_write_5_bits_inputTBE_state_state;
            end else begin
              TBEMemory_15_state_state <= _GEN_2536;
            end
          end else begin
            TBEMemory_15_state_state <= _GEN_2536;
          end
        end else if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_state_state <= io_write_6_bits_inputTBE_state_state;
        end else if (isAlloc_5) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEMemory_15_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_15_state_state <= _GEN_2536;
          end
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_state_state <= 2'h0;
          end else begin
            TBEMemory_15_state_state <= _GEN_2536;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_15_state_state <= _GEN_2536;
          end else if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_state_state <= io_write_5_bits_inputTBE_state_state;
          end else begin
            TBEMemory_15_state_state <= _GEN_2536;
          end
        end else begin
          TBEMemory_15_state_state <= _GEN_2536;
        end
      end else begin
        TBEMemory_15_state_state <= _GEN_3050;
      end
    end else if (_T_243) begin
      if (4'hf == idxUpdate_7[3:0]) begin
        TBEMemory_15_state_state <= 2'h0;
      end else if (isAlloc_6) begin
        if (4'hf == idxAlloc[3:0]) begin
          TBEMemory_15_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_15_state_state <= _GEN_3050;
        end
      end else if (_T_221) begin
        if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_state_state <= 2'h0;
        end else begin
          TBEMemory_15_state_state <= _GEN_3050;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_15_state_state <= _GEN_3050;
        end else if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_15_state_state <= _GEN_3050;
        end
      end else begin
        TBEMemory_15_state_state <= _GEN_3050;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEMemory_15_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_15_state_state <= _GEN_3050;
          end
        end else if (_T_221) begin
          if (4'hf == idxUpdate_6[3:0]) begin
            TBEMemory_15_state_state <= 2'h0;
          end else begin
            TBEMemory_15_state_state <= _GEN_3050;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_15_state_state <= _GEN_3050;
          end else if (4'hf == idxUpdate_6[3:0]) begin
            TBEMemory_15_state_state <= io_write_6_bits_inputTBE_state_state;
          end else begin
            TBEMemory_15_state_state <= _GEN_3050;
          end
        end else begin
          TBEMemory_15_state_state <= _GEN_3050;
        end
      end else if (4'hf == idxUpdate_7[3:0]) begin
        TBEMemory_15_state_state <= io_write_7_bits_inputTBE_state_state;
      end else if (isAlloc_6) begin
        if (4'hf == idxAlloc[3:0]) begin
          TBEMemory_15_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_15_state_state <= _GEN_3050;
        end
      end else if (_T_221) begin
        if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_state_state <= 2'h0;
        end else begin
          TBEMemory_15_state_state <= _GEN_3050;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_15_state_state <= _GEN_3050;
        end else if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_state_state <= io_write_6_bits_inputTBE_state_state;
        end else begin
          TBEMemory_15_state_state <= _GEN_3050;
        end
      end else begin
        TBEMemory_15_state_state <= _GEN_3050;
      end
    end else begin
      TBEMemory_15_state_state <= _GEN_3564;
    end
    if (reset) begin
      TBEMemory_15_way <= 3'h2;
    end else if (isAlloc_7) begin
      if (4'hf == idxAlloc[3:0]) begin
        TBEMemory_15_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'hf == idxAlloc[3:0]) begin
          TBEMemory_15_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEMemory_15_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEMemory_15_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEMemory_15_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEMemory_15_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEMemory_15_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEMemory_15_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEMemory_15_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hf == idxUpdate_0[3:0]) begin
                        TBEMemory_15_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_way <= 3'h2;
                  end else if (isAlloc_0) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEMemory_15_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEMemory_15_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hf == idxUpdate_0[3:0]) begin
                        TBEMemory_15_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (isAlloc_0) begin
                      if (4'hf == idxAlloc[3:0]) begin
                        TBEMemory_15_way <= io_write_0_bits_inputTBE_way;
                      end
                    end else if (_T_89) begin
                      if (4'hf == idxUpdate_0[3:0]) begin
                        TBEMemory_15_way <= 3'h2;
                      end
                    end else if (_T_97) begin
                      if (!(_T_98)) begin
                        if (4'hf == idxUpdate_0[3:0]) begin
                          TBEMemory_15_way <= io_write_0_bits_inputTBE_way;
                        end
                      end
                    end
                  end else if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_way <= io_write_1_bits_inputTBE_way;
                  end else if (isAlloc_0) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEMemory_15_way <= io_write_0_bits_inputTBE_way;
                    end
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEMemory_15_way <= 3'h2;
                    end
                  end else if (_T_97) begin
                    if (!(_T_98)) begin
                      if (4'hf == idxUpdate_0[3:0]) begin
                        TBEMemory_15_way <= io_write_0_bits_inputTBE_way;
                      end
                    end
                  end
                end else begin
                  TBEMemory_15_way <= _GEN_464;
                end
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_way <= 3'h2;
                end else if (isAlloc_1) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEMemory_15_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_15_way <= _GEN_464;
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_way <= 3'h2;
                  end else begin
                    TBEMemory_15_way <= _GEN_464;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_15_way <= _GEN_464;
                  end else if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_15_way <= _GEN_464;
                  end
                end else begin
                  TBEMemory_15_way <= _GEN_464;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (isAlloc_1) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEMemory_15_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_15_way <= _GEN_464;
                    end
                  end else if (_T_111) begin
                    if (4'hf == idxUpdate_1[3:0]) begin
                      TBEMemory_15_way <= 3'h2;
                    end else begin
                      TBEMemory_15_way <= _GEN_464;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      TBEMemory_15_way <= _GEN_464;
                    end else if (4'hf == idxUpdate_1[3:0]) begin
                      TBEMemory_15_way <= io_write_1_bits_inputTBE_way;
                    end else begin
                      TBEMemory_15_way <= _GEN_464;
                    end
                  end else begin
                    TBEMemory_15_way <= _GEN_464;
                  end
                end else if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_way <= io_write_2_bits_inputTBE_way;
                end else if (isAlloc_1) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEMemory_15_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_15_way <= _GEN_464;
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_way <= 3'h2;
                  end else begin
                    TBEMemory_15_way <= _GEN_464;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    TBEMemory_15_way <= _GEN_464;
                  end else if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_way <= io_write_1_bits_inputTBE_way;
                  end else begin
                    TBEMemory_15_way <= _GEN_464;
                  end
                end else begin
                  TBEMemory_15_way <= _GEN_464;
                end
              end else begin
                TBEMemory_15_way <= _GEN_978;
              end
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_way <= 3'h2;
              end else if (isAlloc_2) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEMemory_15_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_15_way <= _GEN_978;
                end
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_way <= 3'h2;
                end else begin
                  TBEMemory_15_way <= _GEN_978;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_15_way <= _GEN_978;
                end else if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_15_way <= _GEN_978;
                end
              end else begin
                TBEMemory_15_way <= _GEN_978;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (isAlloc_2) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEMemory_15_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_15_way <= _GEN_978;
                  end
                end else if (_T_133) begin
                  if (4'hf == idxUpdate_2[3:0]) begin
                    TBEMemory_15_way <= 3'h2;
                  end else begin
                    TBEMemory_15_way <= _GEN_978;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    TBEMemory_15_way <= _GEN_978;
                  end else if (4'hf == idxUpdate_2[3:0]) begin
                    TBEMemory_15_way <= io_write_2_bits_inputTBE_way;
                  end else begin
                    TBEMemory_15_way <= _GEN_978;
                  end
                end else begin
                  TBEMemory_15_way <= _GEN_978;
                end
              end else if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_way <= io_write_3_bits_inputTBE_way;
              end else if (isAlloc_2) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEMemory_15_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_15_way <= _GEN_978;
                end
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_way <= 3'h2;
                end else begin
                  TBEMemory_15_way <= _GEN_978;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  TBEMemory_15_way <= _GEN_978;
                end else if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_way <= io_write_2_bits_inputTBE_way;
                end else begin
                  TBEMemory_15_way <= _GEN_978;
                end
              end else begin
                TBEMemory_15_way <= _GEN_978;
              end
            end else begin
              TBEMemory_15_way <= _GEN_1492;
            end
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_way <= 3'h2;
            end else if (isAlloc_3) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEMemory_15_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_15_way <= _GEN_1492;
              end
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_way <= 3'h2;
              end else begin
                TBEMemory_15_way <= _GEN_1492;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_15_way <= _GEN_1492;
              end else if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_15_way <= _GEN_1492;
              end
            end else begin
              TBEMemory_15_way <= _GEN_1492;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (isAlloc_3) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEMemory_15_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_15_way <= _GEN_1492;
                end
              end else if (_T_155) begin
                if (4'hf == idxUpdate_3[3:0]) begin
                  TBEMemory_15_way <= 3'h2;
                end else begin
                  TBEMemory_15_way <= _GEN_1492;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  TBEMemory_15_way <= _GEN_1492;
                end else if (4'hf == idxUpdate_3[3:0]) begin
                  TBEMemory_15_way <= io_write_3_bits_inputTBE_way;
                end else begin
                  TBEMemory_15_way <= _GEN_1492;
                end
              end else begin
                TBEMemory_15_way <= _GEN_1492;
              end
            end else if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_way <= io_write_4_bits_inputTBE_way;
            end else if (isAlloc_3) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEMemory_15_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_15_way <= _GEN_1492;
              end
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_way <= 3'h2;
              end else begin
                TBEMemory_15_way <= _GEN_1492;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                TBEMemory_15_way <= _GEN_1492;
              end else if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_way <= io_write_3_bits_inputTBE_way;
              end else begin
                TBEMemory_15_way <= _GEN_1492;
              end
            end else begin
              TBEMemory_15_way <= _GEN_1492;
            end
          end else begin
            TBEMemory_15_way <= _GEN_2006;
          end
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_way <= 3'h2;
          end else if (isAlloc_4) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEMemory_15_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_15_way <= _GEN_2006;
            end
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_way <= 3'h2;
            end else begin
              TBEMemory_15_way <= _GEN_2006;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_15_way <= _GEN_2006;
            end else if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_15_way <= _GEN_2006;
            end
          end else begin
            TBEMemory_15_way <= _GEN_2006;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (isAlloc_4) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEMemory_15_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_15_way <= _GEN_2006;
              end
            end else if (_T_177) begin
              if (4'hf == idxUpdate_4[3:0]) begin
                TBEMemory_15_way <= 3'h2;
              end else begin
                TBEMemory_15_way <= _GEN_2006;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                TBEMemory_15_way <= _GEN_2006;
              end else if (4'hf == idxUpdate_4[3:0]) begin
                TBEMemory_15_way <= io_write_4_bits_inputTBE_way;
              end else begin
                TBEMemory_15_way <= _GEN_2006;
              end
            end else begin
              TBEMemory_15_way <= _GEN_2006;
            end
          end else if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_way <= io_write_5_bits_inputTBE_way;
          end else if (isAlloc_4) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEMemory_15_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_15_way <= _GEN_2006;
            end
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_way <= 3'h2;
            end else begin
              TBEMemory_15_way <= _GEN_2006;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              TBEMemory_15_way <= _GEN_2006;
            end else if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_way <= io_write_4_bits_inputTBE_way;
            end else begin
              TBEMemory_15_way <= _GEN_2006;
            end
          end else begin
            TBEMemory_15_way <= _GEN_2006;
          end
        end else begin
          TBEMemory_15_way <= _GEN_2520;
        end
      end else if (_T_221) begin
        if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_way <= 3'h2;
        end else if (isAlloc_5) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEMemory_15_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_15_way <= _GEN_2520;
          end
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_way <= 3'h2;
          end else begin
            TBEMemory_15_way <= _GEN_2520;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_15_way <= _GEN_2520;
          end else if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_15_way <= _GEN_2520;
          end
        end else begin
          TBEMemory_15_way <= _GEN_2520;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (isAlloc_5) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEMemory_15_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_15_way <= _GEN_2520;
            end
          end else if (_T_199) begin
            if (4'hf == idxUpdate_5[3:0]) begin
              TBEMemory_15_way <= 3'h2;
            end else begin
              TBEMemory_15_way <= _GEN_2520;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              TBEMemory_15_way <= _GEN_2520;
            end else if (4'hf == idxUpdate_5[3:0]) begin
              TBEMemory_15_way <= io_write_5_bits_inputTBE_way;
            end else begin
              TBEMemory_15_way <= _GEN_2520;
            end
          end else begin
            TBEMemory_15_way <= _GEN_2520;
          end
        end else if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_way <= io_write_6_bits_inputTBE_way;
        end else if (isAlloc_5) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEMemory_15_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_15_way <= _GEN_2520;
          end
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_way <= 3'h2;
          end else begin
            TBEMemory_15_way <= _GEN_2520;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            TBEMemory_15_way <= _GEN_2520;
          end else if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_way <= io_write_5_bits_inputTBE_way;
          end else begin
            TBEMemory_15_way <= _GEN_2520;
          end
        end else begin
          TBEMemory_15_way <= _GEN_2520;
        end
      end else begin
        TBEMemory_15_way <= _GEN_3034;
      end
    end else if (_T_243) begin
      if (4'hf == idxUpdate_7[3:0]) begin
        TBEMemory_15_way <= 3'h2;
      end else if (isAlloc_6) begin
        if (4'hf == idxAlloc[3:0]) begin
          TBEMemory_15_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_15_way <= _GEN_3034;
        end
      end else if (_T_221) begin
        if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_way <= 3'h2;
        end else begin
          TBEMemory_15_way <= _GEN_3034;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_15_way <= _GEN_3034;
        end else if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_15_way <= _GEN_3034;
        end
      end else begin
        TBEMemory_15_way <= _GEN_3034;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (isAlloc_6) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEMemory_15_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_15_way <= _GEN_3034;
          end
        end else if (_T_221) begin
          if (4'hf == idxUpdate_6[3:0]) begin
            TBEMemory_15_way <= 3'h2;
          end else begin
            TBEMemory_15_way <= _GEN_3034;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            TBEMemory_15_way <= _GEN_3034;
          end else if (4'hf == idxUpdate_6[3:0]) begin
            TBEMemory_15_way <= io_write_6_bits_inputTBE_way;
          end else begin
            TBEMemory_15_way <= _GEN_3034;
          end
        end else begin
          TBEMemory_15_way <= _GEN_3034;
        end
      end else if (4'hf == idxUpdate_7[3:0]) begin
        TBEMemory_15_way <= io_write_7_bits_inputTBE_way;
      end else if (isAlloc_6) begin
        if (4'hf == idxAlloc[3:0]) begin
          TBEMemory_15_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_15_way <= _GEN_3034;
        end
      end else if (_T_221) begin
        if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_way <= 3'h2;
        end else begin
          TBEMemory_15_way <= _GEN_3034;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          TBEMemory_15_way <= _GEN_3034;
        end else if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_way <= io_write_6_bits_inputTBE_way;
        end else begin
          TBEMemory_15_way <= _GEN_3034;
        end
      end else begin
        TBEMemory_15_way <= _GEN_3034;
      end
    end else begin
      TBEMemory_15_way <= _GEN_3548;
    end
    if (reset) begin
      TBEMemory_15_fields_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'hf == idxAlloc[3:0]) begin
        TBEMemory_15_fields_0 <= io_write_7_bits_inputTBE_fields_0;
      end else if (isAlloc_6) begin
        if (4'hf == idxAlloc[3:0]) begin
          TBEMemory_15_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else if (isAlloc_5) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEMemory_15_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else if (isAlloc_4) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEMemory_15_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else if (isAlloc_3) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEMemory_15_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else if (isAlloc_2) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEMemory_15_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else if (isAlloc_1) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEMemory_15_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else if (isAlloc_0) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEMemory_15_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEMemory_15_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'hf == idxUpdate_0[3:0]) begin
                        TBEMemory_15_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_fields_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEMemory_15_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEMemory_15_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'hf == idxUpdate_0[3:0]) begin
                        TBEMemory_15_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'hf == idxUpdate_1[3:0]) begin
                      TBEMemory_15_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else if (isAlloc_0) begin
                      if (4'hf == idxAlloc[3:0]) begin
                        TBEMemory_15_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end else if (_T_89) begin
                      if (4'hf == idxUpdate_0[3:0]) begin
                        TBEMemory_15_fields_0 <= 32'h0;
                      end
                    end else if (_T_97) begin
                      if (_T_98) begin
                        if (4'hf == idxUpdate_0[3:0]) begin
                          TBEMemory_15_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                        end
                      end
                    end
                  end else if (isAlloc_0) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEMemory_15_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                    end
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEMemory_15_fields_0 <= 32'h0;
                    end
                  end else if (_T_97) begin
                    if (_T_98) begin
                      if (4'hf == idxUpdate_0[3:0]) begin
                        TBEMemory_15_fields_0 <= io_write_0_bits_inputTBE_fields_0;
                      end
                    end
                  end
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_448;
                end
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_fields_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEMemory_15_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_448;
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_448;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'hf == idxUpdate_1[3:0]) begin
                      TBEMemory_15_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_15_fields_0 <= _GEN_448;
                    end
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_448;
                  end
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_448;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'hf == idxUpdate_2[3:0]) begin
                    TBEMemory_15_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else if (isAlloc_1) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEMemory_15_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_15_fields_0 <= _GEN_448;
                    end
                  end else if (_T_111) begin
                    if (4'hf == idxUpdate_1[3:0]) begin
                      TBEMemory_15_fields_0 <= 32'h0;
                    end else begin
                      TBEMemory_15_fields_0 <= _GEN_448;
                    end
                  end else if (_T_119) begin
                    if (_T_120) begin
                      if (4'hf == idxUpdate_1[3:0]) begin
                        TBEMemory_15_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                      end else begin
                        TBEMemory_15_fields_0 <= _GEN_448;
                      end
                    end else begin
                      TBEMemory_15_fields_0 <= _GEN_448;
                    end
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_448;
                  end
                end else if (isAlloc_1) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEMemory_15_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_448;
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEMemory_15_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_448;
                  end
                end else if (_T_119) begin
                  if (_T_120) begin
                    if (4'hf == idxUpdate_1[3:0]) begin
                      TBEMemory_15_fields_0 <= io_write_1_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_15_fields_0 <= _GEN_448;
                    end
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_448;
                  end
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_448;
                end
              end else begin
                TBEMemory_15_fields_0 <= _GEN_962;
              end
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_fields_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEMemory_15_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_962;
                end
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_962;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'hf == idxUpdate_2[3:0]) begin
                    TBEMemory_15_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_962;
                  end
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_962;
                end
              end else begin
                TBEMemory_15_fields_0 <= _GEN_962;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'hf == idxUpdate_3[3:0]) begin
                  TBEMemory_15_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else if (isAlloc_2) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEMemory_15_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_962;
                  end
                end else if (_T_133) begin
                  if (4'hf == idxUpdate_2[3:0]) begin
                    TBEMemory_15_fields_0 <= 32'h0;
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_962;
                  end
                end else if (_T_141) begin
                  if (_T_142) begin
                    if (4'hf == idxUpdate_2[3:0]) begin
                      TBEMemory_15_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                    end else begin
                      TBEMemory_15_fields_0 <= _GEN_962;
                    end
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_962;
                  end
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_962;
                end
              end else if (isAlloc_2) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEMemory_15_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_962;
                end
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEMemory_15_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_962;
                end
              end else if (_T_141) begin
                if (_T_142) begin
                  if (4'hf == idxUpdate_2[3:0]) begin
                    TBEMemory_15_fields_0 <= io_write_2_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_962;
                  end
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_962;
                end
              end else begin
                TBEMemory_15_fields_0 <= _GEN_962;
              end
            end else begin
              TBEMemory_15_fields_0 <= _GEN_1476;
            end
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_fields_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEMemory_15_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_15_fields_0 <= _GEN_1476;
              end
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_fields_0 <= 32'h0;
              end else begin
                TBEMemory_15_fields_0 <= _GEN_1476;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'hf == idxUpdate_3[3:0]) begin
                  TBEMemory_15_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_1476;
                end
              end else begin
                TBEMemory_15_fields_0 <= _GEN_1476;
              end
            end else begin
              TBEMemory_15_fields_0 <= _GEN_1476;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'hf == idxUpdate_4[3:0]) begin
                TBEMemory_15_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else if (isAlloc_3) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEMemory_15_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_1476;
                end
              end else if (_T_155) begin
                if (4'hf == idxUpdate_3[3:0]) begin
                  TBEMemory_15_fields_0 <= 32'h0;
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_1476;
                end
              end else if (_T_163) begin
                if (_T_164) begin
                  if (4'hf == idxUpdate_3[3:0]) begin
                    TBEMemory_15_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                  end else begin
                    TBEMemory_15_fields_0 <= _GEN_1476;
                  end
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_1476;
                end
              end else begin
                TBEMemory_15_fields_0 <= _GEN_1476;
              end
            end else if (isAlloc_3) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEMemory_15_fields_0 <= io_write_3_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_15_fields_0 <= _GEN_1476;
              end
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEMemory_15_fields_0 <= 32'h0;
              end else begin
                TBEMemory_15_fields_0 <= _GEN_1476;
              end
            end else if (_T_163) begin
              if (_T_164) begin
                if (4'hf == idxUpdate_3[3:0]) begin
                  TBEMemory_15_fields_0 <= io_write_3_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_1476;
                end
              end else begin
                TBEMemory_15_fields_0 <= _GEN_1476;
              end
            end else begin
              TBEMemory_15_fields_0 <= _GEN_1476;
            end
          end else begin
            TBEMemory_15_fields_0 <= _GEN_1990;
          end
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_fields_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEMemory_15_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_15_fields_0 <= _GEN_1990;
            end
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_fields_0 <= 32'h0;
            end else begin
              TBEMemory_15_fields_0 <= _GEN_1990;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'hf == idxUpdate_4[3:0]) begin
                TBEMemory_15_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_15_fields_0 <= _GEN_1990;
              end
            end else begin
              TBEMemory_15_fields_0 <= _GEN_1990;
            end
          end else begin
            TBEMemory_15_fields_0 <= _GEN_1990;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'hf == idxUpdate_5[3:0]) begin
              TBEMemory_15_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else if (isAlloc_4) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEMemory_15_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_15_fields_0 <= _GEN_1990;
              end
            end else if (_T_177) begin
              if (4'hf == idxUpdate_4[3:0]) begin
                TBEMemory_15_fields_0 <= 32'h0;
              end else begin
                TBEMemory_15_fields_0 <= _GEN_1990;
              end
            end else if (_T_185) begin
              if (_T_186) begin
                if (4'hf == idxUpdate_4[3:0]) begin
                  TBEMemory_15_fields_0 <= io_write_4_bits_inputTBE_fields_0;
                end else begin
                  TBEMemory_15_fields_0 <= _GEN_1990;
                end
              end else begin
                TBEMemory_15_fields_0 <= _GEN_1990;
              end
            end else begin
              TBEMemory_15_fields_0 <= _GEN_1990;
            end
          end else if (isAlloc_4) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEMemory_15_fields_0 <= io_write_4_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_15_fields_0 <= _GEN_1990;
            end
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEMemory_15_fields_0 <= 32'h0;
            end else begin
              TBEMemory_15_fields_0 <= _GEN_1990;
            end
          end else if (_T_185) begin
            if (_T_186) begin
              if (4'hf == idxUpdate_4[3:0]) begin
                TBEMemory_15_fields_0 <= io_write_4_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_15_fields_0 <= _GEN_1990;
              end
            end else begin
              TBEMemory_15_fields_0 <= _GEN_1990;
            end
          end else begin
            TBEMemory_15_fields_0 <= _GEN_1990;
          end
        end else begin
          TBEMemory_15_fields_0 <= _GEN_2504;
        end
      end else if (_T_221) begin
        if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_fields_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEMemory_15_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_15_fields_0 <= _GEN_2504;
          end
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_fields_0 <= 32'h0;
          end else begin
            TBEMemory_15_fields_0 <= _GEN_2504;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'hf == idxUpdate_5[3:0]) begin
              TBEMemory_15_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_15_fields_0 <= _GEN_2504;
            end
          end else begin
            TBEMemory_15_fields_0 <= _GEN_2504;
          end
        end else begin
          TBEMemory_15_fields_0 <= _GEN_2504;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'hf == idxUpdate_6[3:0]) begin
            TBEMemory_15_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else if (isAlloc_5) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEMemory_15_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_15_fields_0 <= _GEN_2504;
            end
          end else if (_T_199) begin
            if (4'hf == idxUpdate_5[3:0]) begin
              TBEMemory_15_fields_0 <= 32'h0;
            end else begin
              TBEMemory_15_fields_0 <= _GEN_2504;
            end
          end else if (_T_207) begin
            if (_T_208) begin
              if (4'hf == idxUpdate_5[3:0]) begin
                TBEMemory_15_fields_0 <= io_write_5_bits_inputTBE_fields_0;
              end else begin
                TBEMemory_15_fields_0 <= _GEN_2504;
              end
            end else begin
              TBEMemory_15_fields_0 <= _GEN_2504;
            end
          end else begin
            TBEMemory_15_fields_0 <= _GEN_2504;
          end
        end else if (isAlloc_5) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEMemory_15_fields_0 <= io_write_5_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_15_fields_0 <= _GEN_2504;
          end
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEMemory_15_fields_0 <= 32'h0;
          end else begin
            TBEMemory_15_fields_0 <= _GEN_2504;
          end
        end else if (_T_207) begin
          if (_T_208) begin
            if (4'hf == idxUpdate_5[3:0]) begin
              TBEMemory_15_fields_0 <= io_write_5_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_15_fields_0 <= _GEN_2504;
            end
          end else begin
            TBEMemory_15_fields_0 <= _GEN_2504;
          end
        end else begin
          TBEMemory_15_fields_0 <= _GEN_2504;
        end
      end else begin
        TBEMemory_15_fields_0 <= _GEN_3018;
      end
    end else if (_T_243) begin
      if (4'hf == idxUpdate_7[3:0]) begin
        TBEMemory_15_fields_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'hf == idxAlloc[3:0]) begin
          TBEMemory_15_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_15_fields_0 <= _GEN_3018;
        end
      end else if (_T_221) begin
        if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_fields_0 <= 32'h0;
        end else begin
          TBEMemory_15_fields_0 <= _GEN_3018;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'hf == idxUpdate_6[3:0]) begin
            TBEMemory_15_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_15_fields_0 <= _GEN_3018;
          end
        end else begin
          TBEMemory_15_fields_0 <= _GEN_3018;
        end
      end else begin
        TBEMemory_15_fields_0 <= _GEN_3018;
      end
    end else if (_T_251) begin
      if (_T_252) begin
        if (4'hf == idxUpdate_7[3:0]) begin
          TBEMemory_15_fields_0 <= io_write_7_bits_inputTBE_fields_0;
        end else if (isAlloc_6) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEMemory_15_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_15_fields_0 <= _GEN_3018;
          end
        end else if (_T_221) begin
          if (4'hf == idxUpdate_6[3:0]) begin
            TBEMemory_15_fields_0 <= 32'h0;
          end else begin
            TBEMemory_15_fields_0 <= _GEN_3018;
          end
        end else if (_T_229) begin
          if (_T_230) begin
            if (4'hf == idxUpdate_6[3:0]) begin
              TBEMemory_15_fields_0 <= io_write_6_bits_inputTBE_fields_0;
            end else begin
              TBEMemory_15_fields_0 <= _GEN_3018;
            end
          end else begin
            TBEMemory_15_fields_0 <= _GEN_3018;
          end
        end else begin
          TBEMemory_15_fields_0 <= _GEN_3018;
        end
      end else if (isAlloc_6) begin
        if (4'hf == idxAlloc[3:0]) begin
          TBEMemory_15_fields_0 <= io_write_6_bits_inputTBE_fields_0;
        end else begin
          TBEMemory_15_fields_0 <= _GEN_3018;
        end
      end else if (_T_221) begin
        if (4'hf == idxUpdate_6[3:0]) begin
          TBEMemory_15_fields_0 <= 32'h0;
        end else begin
          TBEMemory_15_fields_0 <= _GEN_3018;
        end
      end else if (_T_229) begin
        if (_T_230) begin
          if (4'hf == idxUpdate_6[3:0]) begin
            TBEMemory_15_fields_0 <= io_write_6_bits_inputTBE_fields_0;
          end else begin
            TBEMemory_15_fields_0 <= _GEN_3018;
          end
        end else begin
          TBEMemory_15_fields_0 <= _GEN_3018;
        end
      end else begin
        TBEMemory_15_fields_0 <= _GEN_3018;
      end
    end else begin
      TBEMemory_15_fields_0 <= _GEN_3532;
    end
    if (reset) begin
      TBEValid_0 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_0 <= _GEN_3662;
    end else if (_T_243) begin
      if (4'h0 == idxUpdate_7[3:0]) begin
        TBEValid_0 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_0 <= _GEN_3148;
      end else if (_T_221) begin
        if (4'h0 == idxUpdate_6[3:0]) begin
          TBEValid_0 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_0 <= _GEN_2634;
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEValid_0 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_0 <= _GEN_2120;
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEValid_0 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_0 <= _GEN_1606;
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEValid_0 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_0 <= _GEN_1092;
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEValid_0 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_0 <= _GEN_578;
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEValid_0 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_0 <= _GEN_64;
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEValid_0 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_0 <= _GEN_64;
                end else if (_T_89) begin
                  if (4'h0 == idxUpdate_0[3:0]) begin
                    TBEValid_0 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_0 <= _GEN_578;
              end else if (_T_111) begin
                if (4'h0 == idxUpdate_1[3:0]) begin
                  TBEValid_0 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_0 <= _GEN_64;
                end else if (_T_89) begin
                  if (4'h0 == idxUpdate_0[3:0]) begin
                    TBEValid_0 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_0 <= _GEN_64;
              end else if (_T_89) begin
                if (4'h0 == idxUpdate_0[3:0]) begin
                  TBEValid_0 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_0 <= _GEN_1092;
            end else if (_T_133) begin
              if (4'h0 == idxUpdate_2[3:0]) begin
                TBEValid_0 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_0 <= _GEN_578;
              end else if (_T_111) begin
                if (4'h0 == idxUpdate_1[3:0]) begin
                  TBEValid_0 <= 1'h0;
                end else begin
                  TBEValid_0 <= _GEN_497;
                end
              end else begin
                TBEValid_0 <= _GEN_497;
              end
            end else if (isAlloc_1) begin
              TBEValid_0 <= _GEN_578;
            end else if (_T_111) begin
              if (4'h0 == idxUpdate_1[3:0]) begin
                TBEValid_0 <= 1'h0;
              end else begin
                TBEValid_0 <= _GEN_497;
              end
            end else begin
              TBEValid_0 <= _GEN_497;
            end
          end else if (isAlloc_3) begin
            TBEValid_0 <= _GEN_1606;
          end else if (_T_155) begin
            if (4'h0 == idxUpdate_3[3:0]) begin
              TBEValid_0 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_0 <= _GEN_1092;
            end else if (_T_133) begin
              if (4'h0 == idxUpdate_2[3:0]) begin
                TBEValid_0 <= 1'h0;
              end else begin
                TBEValid_0 <= _GEN_1011;
              end
            end else begin
              TBEValid_0 <= _GEN_1011;
            end
          end else if (isAlloc_2) begin
            TBEValid_0 <= _GEN_1092;
          end else if (_T_133) begin
            if (4'h0 == idxUpdate_2[3:0]) begin
              TBEValid_0 <= 1'h0;
            end else begin
              TBEValid_0 <= _GEN_1011;
            end
          end else begin
            TBEValid_0 <= _GEN_1011;
          end
        end else if (isAlloc_4) begin
          TBEValid_0 <= _GEN_2120;
        end else if (_T_177) begin
          if (4'h0 == idxUpdate_4[3:0]) begin
            TBEValid_0 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_0 <= _GEN_1606;
          end else if (_T_155) begin
            if (4'h0 == idxUpdate_3[3:0]) begin
              TBEValid_0 <= 1'h0;
            end else begin
              TBEValid_0 <= _GEN_1525;
            end
          end else begin
            TBEValid_0 <= _GEN_1525;
          end
        end else if (isAlloc_3) begin
          TBEValid_0 <= _GEN_1606;
        end else if (_T_155) begin
          if (4'h0 == idxUpdate_3[3:0]) begin
            TBEValid_0 <= 1'h0;
          end else begin
            TBEValid_0 <= _GEN_1525;
          end
        end else begin
          TBEValid_0 <= _GEN_1525;
        end
      end else if (isAlloc_5) begin
        TBEValid_0 <= _GEN_2634;
      end else if (_T_199) begin
        if (4'h0 == idxUpdate_5[3:0]) begin
          TBEValid_0 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_0 <= _GEN_2120;
        end else if (_T_177) begin
          if (4'h0 == idxUpdate_4[3:0]) begin
            TBEValid_0 <= 1'h0;
          end else begin
            TBEValid_0 <= _GEN_2039;
          end
        end else begin
          TBEValid_0 <= _GEN_2039;
        end
      end else if (isAlloc_4) begin
        TBEValid_0 <= _GEN_2120;
      end else if (_T_177) begin
        if (4'h0 == idxUpdate_4[3:0]) begin
          TBEValid_0 <= 1'h0;
        end else begin
          TBEValid_0 <= _GEN_2039;
        end
      end else begin
        TBEValid_0 <= _GEN_2039;
      end
    end else if (isAlloc_6) begin
      TBEValid_0 <= _GEN_3148;
    end else if (_T_221) begin
      if (4'h0 == idxUpdate_6[3:0]) begin
        TBEValid_0 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_0 <= _GEN_2634;
      end else if (_T_199) begin
        if (4'h0 == idxUpdate_5[3:0]) begin
          TBEValid_0 <= 1'h0;
        end else begin
          TBEValid_0 <= _GEN_2553;
        end
      end else begin
        TBEValid_0 <= _GEN_2553;
      end
    end else if (isAlloc_5) begin
      TBEValid_0 <= _GEN_2634;
    end else if (_T_199) begin
      if (4'h0 == idxUpdate_5[3:0]) begin
        TBEValid_0 <= 1'h0;
      end else begin
        TBEValid_0 <= _GEN_2553;
      end
    end else begin
      TBEValid_0 <= _GEN_2553;
    end
    if (reset) begin
      TBEValid_1 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_1 <= _GEN_3663;
    end else if (_T_243) begin
      if (4'h1 == idxUpdate_7[3:0]) begin
        TBEValid_1 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_1 <= _GEN_3149;
      end else if (_T_221) begin
        if (4'h1 == idxUpdate_6[3:0]) begin
          TBEValid_1 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_1 <= _GEN_2635;
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEValid_1 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_1 <= _GEN_2121;
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEValid_1 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_1 <= _GEN_1607;
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEValid_1 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_1 <= _GEN_1093;
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEValid_1 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_1 <= _GEN_579;
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEValid_1 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_1 <= _GEN_65;
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEValid_1 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_1 <= _GEN_65;
                end else if (_T_89) begin
                  if (4'h1 == idxUpdate_0[3:0]) begin
                    TBEValid_1 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_1 <= _GEN_579;
              end else if (_T_111) begin
                if (4'h1 == idxUpdate_1[3:0]) begin
                  TBEValid_1 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_1 <= _GEN_65;
                end else if (_T_89) begin
                  if (4'h1 == idxUpdate_0[3:0]) begin
                    TBEValid_1 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_1 <= _GEN_65;
              end else if (_T_89) begin
                if (4'h1 == idxUpdate_0[3:0]) begin
                  TBEValid_1 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_1 <= _GEN_1093;
            end else if (_T_133) begin
              if (4'h1 == idxUpdate_2[3:0]) begin
                TBEValid_1 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_1 <= _GEN_579;
              end else if (_T_111) begin
                if (4'h1 == idxUpdate_1[3:0]) begin
                  TBEValid_1 <= 1'h0;
                end else begin
                  TBEValid_1 <= _GEN_498;
                end
              end else begin
                TBEValid_1 <= _GEN_498;
              end
            end else if (isAlloc_1) begin
              TBEValid_1 <= _GEN_579;
            end else if (_T_111) begin
              if (4'h1 == idxUpdate_1[3:0]) begin
                TBEValid_1 <= 1'h0;
              end else begin
                TBEValid_1 <= _GEN_498;
              end
            end else begin
              TBEValid_1 <= _GEN_498;
            end
          end else if (isAlloc_3) begin
            TBEValid_1 <= _GEN_1607;
          end else if (_T_155) begin
            if (4'h1 == idxUpdate_3[3:0]) begin
              TBEValid_1 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_1 <= _GEN_1093;
            end else if (_T_133) begin
              if (4'h1 == idxUpdate_2[3:0]) begin
                TBEValid_1 <= 1'h0;
              end else begin
                TBEValid_1 <= _GEN_1012;
              end
            end else begin
              TBEValid_1 <= _GEN_1012;
            end
          end else if (isAlloc_2) begin
            TBEValid_1 <= _GEN_1093;
          end else if (_T_133) begin
            if (4'h1 == idxUpdate_2[3:0]) begin
              TBEValid_1 <= 1'h0;
            end else begin
              TBEValid_1 <= _GEN_1012;
            end
          end else begin
            TBEValid_1 <= _GEN_1012;
          end
        end else if (isAlloc_4) begin
          TBEValid_1 <= _GEN_2121;
        end else if (_T_177) begin
          if (4'h1 == idxUpdate_4[3:0]) begin
            TBEValid_1 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_1 <= _GEN_1607;
          end else if (_T_155) begin
            if (4'h1 == idxUpdate_3[3:0]) begin
              TBEValid_1 <= 1'h0;
            end else begin
              TBEValid_1 <= _GEN_1526;
            end
          end else begin
            TBEValid_1 <= _GEN_1526;
          end
        end else if (isAlloc_3) begin
          TBEValid_1 <= _GEN_1607;
        end else if (_T_155) begin
          if (4'h1 == idxUpdate_3[3:0]) begin
            TBEValid_1 <= 1'h0;
          end else begin
            TBEValid_1 <= _GEN_1526;
          end
        end else begin
          TBEValid_1 <= _GEN_1526;
        end
      end else if (isAlloc_5) begin
        TBEValid_1 <= _GEN_2635;
      end else if (_T_199) begin
        if (4'h1 == idxUpdate_5[3:0]) begin
          TBEValid_1 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_1 <= _GEN_2121;
        end else if (_T_177) begin
          if (4'h1 == idxUpdate_4[3:0]) begin
            TBEValid_1 <= 1'h0;
          end else begin
            TBEValid_1 <= _GEN_2040;
          end
        end else begin
          TBEValid_1 <= _GEN_2040;
        end
      end else if (isAlloc_4) begin
        TBEValid_1 <= _GEN_2121;
      end else if (_T_177) begin
        if (4'h1 == idxUpdate_4[3:0]) begin
          TBEValid_1 <= 1'h0;
        end else begin
          TBEValid_1 <= _GEN_2040;
        end
      end else begin
        TBEValid_1 <= _GEN_2040;
      end
    end else if (isAlloc_6) begin
      TBEValid_1 <= _GEN_3149;
    end else if (_T_221) begin
      if (4'h1 == idxUpdate_6[3:0]) begin
        TBEValid_1 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_1 <= _GEN_2635;
      end else if (_T_199) begin
        if (4'h1 == idxUpdate_5[3:0]) begin
          TBEValid_1 <= 1'h0;
        end else begin
          TBEValid_1 <= _GEN_2554;
        end
      end else begin
        TBEValid_1 <= _GEN_2554;
      end
    end else if (isAlloc_5) begin
      TBEValid_1 <= _GEN_2635;
    end else if (_T_199) begin
      if (4'h1 == idxUpdate_5[3:0]) begin
        TBEValid_1 <= 1'h0;
      end else begin
        TBEValid_1 <= _GEN_2554;
      end
    end else begin
      TBEValid_1 <= _GEN_2554;
    end
    if (reset) begin
      TBEValid_2 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_2 <= _GEN_3664;
    end else if (_T_243) begin
      if (4'h2 == idxUpdate_7[3:0]) begin
        TBEValid_2 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_2 <= _GEN_3150;
      end else if (_T_221) begin
        if (4'h2 == idxUpdate_6[3:0]) begin
          TBEValid_2 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_2 <= _GEN_2636;
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEValid_2 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_2 <= _GEN_2122;
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEValid_2 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_2 <= _GEN_1608;
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEValid_2 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_2 <= _GEN_1094;
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEValid_2 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_2 <= _GEN_580;
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEValid_2 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_2 <= _GEN_66;
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEValid_2 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_2 <= _GEN_66;
                end else if (_T_89) begin
                  if (4'h2 == idxUpdate_0[3:0]) begin
                    TBEValid_2 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_2 <= _GEN_580;
              end else if (_T_111) begin
                if (4'h2 == idxUpdate_1[3:0]) begin
                  TBEValid_2 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_2 <= _GEN_66;
                end else if (_T_89) begin
                  if (4'h2 == idxUpdate_0[3:0]) begin
                    TBEValid_2 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_2 <= _GEN_66;
              end else if (_T_89) begin
                if (4'h2 == idxUpdate_0[3:0]) begin
                  TBEValid_2 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_2 <= _GEN_1094;
            end else if (_T_133) begin
              if (4'h2 == idxUpdate_2[3:0]) begin
                TBEValid_2 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_2 <= _GEN_580;
              end else if (_T_111) begin
                if (4'h2 == idxUpdate_1[3:0]) begin
                  TBEValid_2 <= 1'h0;
                end else begin
                  TBEValid_2 <= _GEN_499;
                end
              end else begin
                TBEValid_2 <= _GEN_499;
              end
            end else if (isAlloc_1) begin
              TBEValid_2 <= _GEN_580;
            end else if (_T_111) begin
              if (4'h2 == idxUpdate_1[3:0]) begin
                TBEValid_2 <= 1'h0;
              end else begin
                TBEValid_2 <= _GEN_499;
              end
            end else begin
              TBEValid_2 <= _GEN_499;
            end
          end else if (isAlloc_3) begin
            TBEValid_2 <= _GEN_1608;
          end else if (_T_155) begin
            if (4'h2 == idxUpdate_3[3:0]) begin
              TBEValid_2 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_2 <= _GEN_1094;
            end else if (_T_133) begin
              if (4'h2 == idxUpdate_2[3:0]) begin
                TBEValid_2 <= 1'h0;
              end else begin
                TBEValid_2 <= _GEN_1013;
              end
            end else begin
              TBEValid_2 <= _GEN_1013;
            end
          end else if (isAlloc_2) begin
            TBEValid_2 <= _GEN_1094;
          end else if (_T_133) begin
            if (4'h2 == idxUpdate_2[3:0]) begin
              TBEValid_2 <= 1'h0;
            end else begin
              TBEValid_2 <= _GEN_1013;
            end
          end else begin
            TBEValid_2 <= _GEN_1013;
          end
        end else if (isAlloc_4) begin
          TBEValid_2 <= _GEN_2122;
        end else if (_T_177) begin
          if (4'h2 == idxUpdate_4[3:0]) begin
            TBEValid_2 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_2 <= _GEN_1608;
          end else if (_T_155) begin
            if (4'h2 == idxUpdate_3[3:0]) begin
              TBEValid_2 <= 1'h0;
            end else begin
              TBEValid_2 <= _GEN_1527;
            end
          end else begin
            TBEValid_2 <= _GEN_1527;
          end
        end else if (isAlloc_3) begin
          TBEValid_2 <= _GEN_1608;
        end else if (_T_155) begin
          if (4'h2 == idxUpdate_3[3:0]) begin
            TBEValid_2 <= 1'h0;
          end else begin
            TBEValid_2 <= _GEN_1527;
          end
        end else begin
          TBEValid_2 <= _GEN_1527;
        end
      end else if (isAlloc_5) begin
        TBEValid_2 <= _GEN_2636;
      end else if (_T_199) begin
        if (4'h2 == idxUpdate_5[3:0]) begin
          TBEValid_2 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_2 <= _GEN_2122;
        end else if (_T_177) begin
          if (4'h2 == idxUpdate_4[3:0]) begin
            TBEValid_2 <= 1'h0;
          end else begin
            TBEValid_2 <= _GEN_2041;
          end
        end else begin
          TBEValid_2 <= _GEN_2041;
        end
      end else if (isAlloc_4) begin
        TBEValid_2 <= _GEN_2122;
      end else if (_T_177) begin
        if (4'h2 == idxUpdate_4[3:0]) begin
          TBEValid_2 <= 1'h0;
        end else begin
          TBEValid_2 <= _GEN_2041;
        end
      end else begin
        TBEValid_2 <= _GEN_2041;
      end
    end else if (isAlloc_6) begin
      TBEValid_2 <= _GEN_3150;
    end else if (_T_221) begin
      if (4'h2 == idxUpdate_6[3:0]) begin
        TBEValid_2 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_2 <= _GEN_2636;
      end else if (_T_199) begin
        if (4'h2 == idxUpdate_5[3:0]) begin
          TBEValid_2 <= 1'h0;
        end else begin
          TBEValid_2 <= _GEN_2555;
        end
      end else begin
        TBEValid_2 <= _GEN_2555;
      end
    end else if (isAlloc_5) begin
      TBEValid_2 <= _GEN_2636;
    end else if (_T_199) begin
      if (4'h2 == idxUpdate_5[3:0]) begin
        TBEValid_2 <= 1'h0;
      end else begin
        TBEValid_2 <= _GEN_2555;
      end
    end else begin
      TBEValid_2 <= _GEN_2555;
    end
    if (reset) begin
      TBEValid_3 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_3 <= _GEN_3665;
    end else if (_T_243) begin
      if (4'h3 == idxUpdate_7[3:0]) begin
        TBEValid_3 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_3 <= _GEN_3151;
      end else if (_T_221) begin
        if (4'h3 == idxUpdate_6[3:0]) begin
          TBEValid_3 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_3 <= _GEN_2637;
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEValid_3 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_3 <= _GEN_2123;
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEValid_3 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_3 <= _GEN_1609;
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEValid_3 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_3 <= _GEN_1095;
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEValid_3 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_3 <= _GEN_581;
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEValid_3 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_3 <= _GEN_67;
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEValid_3 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_3 <= _GEN_67;
                end else if (_T_89) begin
                  if (4'h3 == idxUpdate_0[3:0]) begin
                    TBEValid_3 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_3 <= _GEN_581;
              end else if (_T_111) begin
                if (4'h3 == idxUpdate_1[3:0]) begin
                  TBEValid_3 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_3 <= _GEN_67;
                end else if (_T_89) begin
                  if (4'h3 == idxUpdate_0[3:0]) begin
                    TBEValid_3 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_3 <= _GEN_67;
              end else if (_T_89) begin
                if (4'h3 == idxUpdate_0[3:0]) begin
                  TBEValid_3 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_3 <= _GEN_1095;
            end else if (_T_133) begin
              if (4'h3 == idxUpdate_2[3:0]) begin
                TBEValid_3 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_3 <= _GEN_581;
              end else if (_T_111) begin
                if (4'h3 == idxUpdate_1[3:0]) begin
                  TBEValid_3 <= 1'h0;
                end else begin
                  TBEValid_3 <= _GEN_500;
                end
              end else begin
                TBEValid_3 <= _GEN_500;
              end
            end else if (isAlloc_1) begin
              TBEValid_3 <= _GEN_581;
            end else if (_T_111) begin
              if (4'h3 == idxUpdate_1[3:0]) begin
                TBEValid_3 <= 1'h0;
              end else begin
                TBEValid_3 <= _GEN_500;
              end
            end else begin
              TBEValid_3 <= _GEN_500;
            end
          end else if (isAlloc_3) begin
            TBEValid_3 <= _GEN_1609;
          end else if (_T_155) begin
            if (4'h3 == idxUpdate_3[3:0]) begin
              TBEValid_3 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_3 <= _GEN_1095;
            end else if (_T_133) begin
              if (4'h3 == idxUpdate_2[3:0]) begin
                TBEValid_3 <= 1'h0;
              end else begin
                TBEValid_3 <= _GEN_1014;
              end
            end else begin
              TBEValid_3 <= _GEN_1014;
            end
          end else if (isAlloc_2) begin
            TBEValid_3 <= _GEN_1095;
          end else if (_T_133) begin
            if (4'h3 == idxUpdate_2[3:0]) begin
              TBEValid_3 <= 1'h0;
            end else begin
              TBEValid_3 <= _GEN_1014;
            end
          end else begin
            TBEValid_3 <= _GEN_1014;
          end
        end else if (isAlloc_4) begin
          TBEValid_3 <= _GEN_2123;
        end else if (_T_177) begin
          if (4'h3 == idxUpdate_4[3:0]) begin
            TBEValid_3 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_3 <= _GEN_1609;
          end else if (_T_155) begin
            if (4'h3 == idxUpdate_3[3:0]) begin
              TBEValid_3 <= 1'h0;
            end else begin
              TBEValid_3 <= _GEN_1528;
            end
          end else begin
            TBEValid_3 <= _GEN_1528;
          end
        end else if (isAlloc_3) begin
          TBEValid_3 <= _GEN_1609;
        end else if (_T_155) begin
          if (4'h3 == idxUpdate_3[3:0]) begin
            TBEValid_3 <= 1'h0;
          end else begin
            TBEValid_3 <= _GEN_1528;
          end
        end else begin
          TBEValid_3 <= _GEN_1528;
        end
      end else if (isAlloc_5) begin
        TBEValid_3 <= _GEN_2637;
      end else if (_T_199) begin
        if (4'h3 == idxUpdate_5[3:0]) begin
          TBEValid_3 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_3 <= _GEN_2123;
        end else if (_T_177) begin
          if (4'h3 == idxUpdate_4[3:0]) begin
            TBEValid_3 <= 1'h0;
          end else begin
            TBEValid_3 <= _GEN_2042;
          end
        end else begin
          TBEValid_3 <= _GEN_2042;
        end
      end else if (isAlloc_4) begin
        TBEValid_3 <= _GEN_2123;
      end else if (_T_177) begin
        if (4'h3 == idxUpdate_4[3:0]) begin
          TBEValid_3 <= 1'h0;
        end else begin
          TBEValid_3 <= _GEN_2042;
        end
      end else begin
        TBEValid_3 <= _GEN_2042;
      end
    end else if (isAlloc_6) begin
      TBEValid_3 <= _GEN_3151;
    end else if (_T_221) begin
      if (4'h3 == idxUpdate_6[3:0]) begin
        TBEValid_3 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_3 <= _GEN_2637;
      end else if (_T_199) begin
        if (4'h3 == idxUpdate_5[3:0]) begin
          TBEValid_3 <= 1'h0;
        end else begin
          TBEValid_3 <= _GEN_2556;
        end
      end else begin
        TBEValid_3 <= _GEN_2556;
      end
    end else if (isAlloc_5) begin
      TBEValid_3 <= _GEN_2637;
    end else if (_T_199) begin
      if (4'h3 == idxUpdate_5[3:0]) begin
        TBEValid_3 <= 1'h0;
      end else begin
        TBEValid_3 <= _GEN_2556;
      end
    end else begin
      TBEValid_3 <= _GEN_2556;
    end
    if (reset) begin
      TBEValid_4 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_4 <= _GEN_3666;
    end else if (_T_243) begin
      if (4'h4 == idxUpdate_7[3:0]) begin
        TBEValid_4 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_4 <= _GEN_3152;
      end else if (_T_221) begin
        if (4'h4 == idxUpdate_6[3:0]) begin
          TBEValid_4 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_4 <= _GEN_2638;
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEValid_4 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_4 <= _GEN_2124;
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEValid_4 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_4 <= _GEN_1610;
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEValid_4 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_4 <= _GEN_1096;
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEValid_4 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_4 <= _GEN_582;
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEValid_4 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_4 <= _GEN_68;
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEValid_4 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_4 <= _GEN_68;
                end else if (_T_89) begin
                  if (4'h4 == idxUpdate_0[3:0]) begin
                    TBEValid_4 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_4 <= _GEN_582;
              end else if (_T_111) begin
                if (4'h4 == idxUpdate_1[3:0]) begin
                  TBEValid_4 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_4 <= _GEN_68;
                end else if (_T_89) begin
                  if (4'h4 == idxUpdate_0[3:0]) begin
                    TBEValid_4 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_4 <= _GEN_68;
              end else if (_T_89) begin
                if (4'h4 == idxUpdate_0[3:0]) begin
                  TBEValid_4 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_4 <= _GEN_1096;
            end else if (_T_133) begin
              if (4'h4 == idxUpdate_2[3:0]) begin
                TBEValid_4 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_4 <= _GEN_582;
              end else if (_T_111) begin
                if (4'h4 == idxUpdate_1[3:0]) begin
                  TBEValid_4 <= 1'h0;
                end else begin
                  TBEValid_4 <= _GEN_501;
                end
              end else begin
                TBEValid_4 <= _GEN_501;
              end
            end else if (isAlloc_1) begin
              TBEValid_4 <= _GEN_582;
            end else if (_T_111) begin
              if (4'h4 == idxUpdate_1[3:0]) begin
                TBEValid_4 <= 1'h0;
              end else begin
                TBEValid_4 <= _GEN_501;
              end
            end else begin
              TBEValid_4 <= _GEN_501;
            end
          end else if (isAlloc_3) begin
            TBEValid_4 <= _GEN_1610;
          end else if (_T_155) begin
            if (4'h4 == idxUpdate_3[3:0]) begin
              TBEValid_4 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_4 <= _GEN_1096;
            end else if (_T_133) begin
              if (4'h4 == idxUpdate_2[3:0]) begin
                TBEValid_4 <= 1'h0;
              end else begin
                TBEValid_4 <= _GEN_1015;
              end
            end else begin
              TBEValid_4 <= _GEN_1015;
            end
          end else if (isAlloc_2) begin
            TBEValid_4 <= _GEN_1096;
          end else if (_T_133) begin
            if (4'h4 == idxUpdate_2[3:0]) begin
              TBEValid_4 <= 1'h0;
            end else begin
              TBEValid_4 <= _GEN_1015;
            end
          end else begin
            TBEValid_4 <= _GEN_1015;
          end
        end else if (isAlloc_4) begin
          TBEValid_4 <= _GEN_2124;
        end else if (_T_177) begin
          if (4'h4 == idxUpdate_4[3:0]) begin
            TBEValid_4 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_4 <= _GEN_1610;
          end else if (_T_155) begin
            if (4'h4 == idxUpdate_3[3:0]) begin
              TBEValid_4 <= 1'h0;
            end else begin
              TBEValid_4 <= _GEN_1529;
            end
          end else begin
            TBEValid_4 <= _GEN_1529;
          end
        end else if (isAlloc_3) begin
          TBEValid_4 <= _GEN_1610;
        end else if (_T_155) begin
          if (4'h4 == idxUpdate_3[3:0]) begin
            TBEValid_4 <= 1'h0;
          end else begin
            TBEValid_4 <= _GEN_1529;
          end
        end else begin
          TBEValid_4 <= _GEN_1529;
        end
      end else if (isAlloc_5) begin
        TBEValid_4 <= _GEN_2638;
      end else if (_T_199) begin
        if (4'h4 == idxUpdate_5[3:0]) begin
          TBEValid_4 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_4 <= _GEN_2124;
        end else if (_T_177) begin
          if (4'h4 == idxUpdate_4[3:0]) begin
            TBEValid_4 <= 1'h0;
          end else begin
            TBEValid_4 <= _GEN_2043;
          end
        end else begin
          TBEValid_4 <= _GEN_2043;
        end
      end else if (isAlloc_4) begin
        TBEValid_4 <= _GEN_2124;
      end else if (_T_177) begin
        if (4'h4 == idxUpdate_4[3:0]) begin
          TBEValid_4 <= 1'h0;
        end else begin
          TBEValid_4 <= _GEN_2043;
        end
      end else begin
        TBEValid_4 <= _GEN_2043;
      end
    end else if (isAlloc_6) begin
      TBEValid_4 <= _GEN_3152;
    end else if (_T_221) begin
      if (4'h4 == idxUpdate_6[3:0]) begin
        TBEValid_4 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_4 <= _GEN_2638;
      end else if (_T_199) begin
        if (4'h4 == idxUpdate_5[3:0]) begin
          TBEValid_4 <= 1'h0;
        end else begin
          TBEValid_4 <= _GEN_2557;
        end
      end else begin
        TBEValid_4 <= _GEN_2557;
      end
    end else if (isAlloc_5) begin
      TBEValid_4 <= _GEN_2638;
    end else if (_T_199) begin
      if (4'h4 == idxUpdate_5[3:0]) begin
        TBEValid_4 <= 1'h0;
      end else begin
        TBEValid_4 <= _GEN_2557;
      end
    end else begin
      TBEValid_4 <= _GEN_2557;
    end
    if (reset) begin
      TBEValid_5 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_5 <= _GEN_3667;
    end else if (_T_243) begin
      if (4'h5 == idxUpdate_7[3:0]) begin
        TBEValid_5 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_5 <= _GEN_3153;
      end else if (_T_221) begin
        if (4'h5 == idxUpdate_6[3:0]) begin
          TBEValid_5 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_5 <= _GEN_2639;
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEValid_5 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_5 <= _GEN_2125;
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEValid_5 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_5 <= _GEN_1611;
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEValid_5 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_5 <= _GEN_1097;
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEValid_5 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_5 <= _GEN_583;
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEValid_5 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_5 <= _GEN_69;
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEValid_5 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_5 <= _GEN_69;
                end else if (_T_89) begin
                  if (4'h5 == idxUpdate_0[3:0]) begin
                    TBEValid_5 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_5 <= _GEN_583;
              end else if (_T_111) begin
                if (4'h5 == idxUpdate_1[3:0]) begin
                  TBEValid_5 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_5 <= _GEN_69;
                end else if (_T_89) begin
                  if (4'h5 == idxUpdate_0[3:0]) begin
                    TBEValid_5 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_5 <= _GEN_69;
              end else if (_T_89) begin
                if (4'h5 == idxUpdate_0[3:0]) begin
                  TBEValid_5 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_5 <= _GEN_1097;
            end else if (_T_133) begin
              if (4'h5 == idxUpdate_2[3:0]) begin
                TBEValid_5 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_5 <= _GEN_583;
              end else if (_T_111) begin
                if (4'h5 == idxUpdate_1[3:0]) begin
                  TBEValid_5 <= 1'h0;
                end else begin
                  TBEValid_5 <= _GEN_502;
                end
              end else begin
                TBEValid_5 <= _GEN_502;
              end
            end else if (isAlloc_1) begin
              TBEValid_5 <= _GEN_583;
            end else if (_T_111) begin
              if (4'h5 == idxUpdate_1[3:0]) begin
                TBEValid_5 <= 1'h0;
              end else begin
                TBEValid_5 <= _GEN_502;
              end
            end else begin
              TBEValid_5 <= _GEN_502;
            end
          end else if (isAlloc_3) begin
            TBEValid_5 <= _GEN_1611;
          end else if (_T_155) begin
            if (4'h5 == idxUpdate_3[3:0]) begin
              TBEValid_5 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_5 <= _GEN_1097;
            end else if (_T_133) begin
              if (4'h5 == idxUpdate_2[3:0]) begin
                TBEValid_5 <= 1'h0;
              end else begin
                TBEValid_5 <= _GEN_1016;
              end
            end else begin
              TBEValid_5 <= _GEN_1016;
            end
          end else if (isAlloc_2) begin
            TBEValid_5 <= _GEN_1097;
          end else if (_T_133) begin
            if (4'h5 == idxUpdate_2[3:0]) begin
              TBEValid_5 <= 1'h0;
            end else begin
              TBEValid_5 <= _GEN_1016;
            end
          end else begin
            TBEValid_5 <= _GEN_1016;
          end
        end else if (isAlloc_4) begin
          TBEValid_5 <= _GEN_2125;
        end else if (_T_177) begin
          if (4'h5 == idxUpdate_4[3:0]) begin
            TBEValid_5 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_5 <= _GEN_1611;
          end else if (_T_155) begin
            if (4'h5 == idxUpdate_3[3:0]) begin
              TBEValid_5 <= 1'h0;
            end else begin
              TBEValid_5 <= _GEN_1530;
            end
          end else begin
            TBEValid_5 <= _GEN_1530;
          end
        end else if (isAlloc_3) begin
          TBEValid_5 <= _GEN_1611;
        end else if (_T_155) begin
          if (4'h5 == idxUpdate_3[3:0]) begin
            TBEValid_5 <= 1'h0;
          end else begin
            TBEValid_5 <= _GEN_1530;
          end
        end else begin
          TBEValid_5 <= _GEN_1530;
        end
      end else if (isAlloc_5) begin
        TBEValid_5 <= _GEN_2639;
      end else if (_T_199) begin
        if (4'h5 == idxUpdate_5[3:0]) begin
          TBEValid_5 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_5 <= _GEN_2125;
        end else if (_T_177) begin
          if (4'h5 == idxUpdate_4[3:0]) begin
            TBEValid_5 <= 1'h0;
          end else begin
            TBEValid_5 <= _GEN_2044;
          end
        end else begin
          TBEValid_5 <= _GEN_2044;
        end
      end else if (isAlloc_4) begin
        TBEValid_5 <= _GEN_2125;
      end else if (_T_177) begin
        if (4'h5 == idxUpdate_4[3:0]) begin
          TBEValid_5 <= 1'h0;
        end else begin
          TBEValid_5 <= _GEN_2044;
        end
      end else begin
        TBEValid_5 <= _GEN_2044;
      end
    end else if (isAlloc_6) begin
      TBEValid_5 <= _GEN_3153;
    end else if (_T_221) begin
      if (4'h5 == idxUpdate_6[3:0]) begin
        TBEValid_5 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_5 <= _GEN_2639;
      end else if (_T_199) begin
        if (4'h5 == idxUpdate_5[3:0]) begin
          TBEValid_5 <= 1'h0;
        end else begin
          TBEValid_5 <= _GEN_2558;
        end
      end else begin
        TBEValid_5 <= _GEN_2558;
      end
    end else if (isAlloc_5) begin
      TBEValid_5 <= _GEN_2639;
    end else if (_T_199) begin
      if (4'h5 == idxUpdate_5[3:0]) begin
        TBEValid_5 <= 1'h0;
      end else begin
        TBEValid_5 <= _GEN_2558;
      end
    end else begin
      TBEValid_5 <= _GEN_2558;
    end
    if (reset) begin
      TBEValid_6 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_6 <= _GEN_3668;
    end else if (_T_243) begin
      if (4'h6 == idxUpdate_7[3:0]) begin
        TBEValid_6 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_6 <= _GEN_3154;
      end else if (_T_221) begin
        if (4'h6 == idxUpdate_6[3:0]) begin
          TBEValid_6 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_6 <= _GEN_2640;
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEValid_6 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_6 <= _GEN_2126;
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEValid_6 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_6 <= _GEN_1612;
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEValid_6 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_6 <= _GEN_1098;
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEValid_6 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_6 <= _GEN_584;
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEValid_6 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_6 <= _GEN_70;
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEValid_6 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_6 <= _GEN_70;
                end else if (_T_89) begin
                  if (4'h6 == idxUpdate_0[3:0]) begin
                    TBEValid_6 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_6 <= _GEN_584;
              end else if (_T_111) begin
                if (4'h6 == idxUpdate_1[3:0]) begin
                  TBEValid_6 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_6 <= _GEN_70;
                end else if (_T_89) begin
                  if (4'h6 == idxUpdate_0[3:0]) begin
                    TBEValid_6 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_6 <= _GEN_70;
              end else if (_T_89) begin
                if (4'h6 == idxUpdate_0[3:0]) begin
                  TBEValid_6 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_6 <= _GEN_1098;
            end else if (_T_133) begin
              if (4'h6 == idxUpdate_2[3:0]) begin
                TBEValid_6 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_6 <= _GEN_584;
              end else if (_T_111) begin
                if (4'h6 == idxUpdate_1[3:0]) begin
                  TBEValid_6 <= 1'h0;
                end else begin
                  TBEValid_6 <= _GEN_503;
                end
              end else begin
                TBEValid_6 <= _GEN_503;
              end
            end else if (isAlloc_1) begin
              TBEValid_6 <= _GEN_584;
            end else if (_T_111) begin
              if (4'h6 == idxUpdate_1[3:0]) begin
                TBEValid_6 <= 1'h0;
              end else begin
                TBEValid_6 <= _GEN_503;
              end
            end else begin
              TBEValid_6 <= _GEN_503;
            end
          end else if (isAlloc_3) begin
            TBEValid_6 <= _GEN_1612;
          end else if (_T_155) begin
            if (4'h6 == idxUpdate_3[3:0]) begin
              TBEValid_6 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_6 <= _GEN_1098;
            end else if (_T_133) begin
              if (4'h6 == idxUpdate_2[3:0]) begin
                TBEValid_6 <= 1'h0;
              end else begin
                TBEValid_6 <= _GEN_1017;
              end
            end else begin
              TBEValid_6 <= _GEN_1017;
            end
          end else if (isAlloc_2) begin
            TBEValid_6 <= _GEN_1098;
          end else if (_T_133) begin
            if (4'h6 == idxUpdate_2[3:0]) begin
              TBEValid_6 <= 1'h0;
            end else begin
              TBEValid_6 <= _GEN_1017;
            end
          end else begin
            TBEValid_6 <= _GEN_1017;
          end
        end else if (isAlloc_4) begin
          TBEValid_6 <= _GEN_2126;
        end else if (_T_177) begin
          if (4'h6 == idxUpdate_4[3:0]) begin
            TBEValid_6 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_6 <= _GEN_1612;
          end else if (_T_155) begin
            if (4'h6 == idxUpdate_3[3:0]) begin
              TBEValid_6 <= 1'h0;
            end else begin
              TBEValid_6 <= _GEN_1531;
            end
          end else begin
            TBEValid_6 <= _GEN_1531;
          end
        end else if (isAlloc_3) begin
          TBEValid_6 <= _GEN_1612;
        end else if (_T_155) begin
          if (4'h6 == idxUpdate_3[3:0]) begin
            TBEValid_6 <= 1'h0;
          end else begin
            TBEValid_6 <= _GEN_1531;
          end
        end else begin
          TBEValid_6 <= _GEN_1531;
        end
      end else if (isAlloc_5) begin
        TBEValid_6 <= _GEN_2640;
      end else if (_T_199) begin
        if (4'h6 == idxUpdate_5[3:0]) begin
          TBEValid_6 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_6 <= _GEN_2126;
        end else if (_T_177) begin
          if (4'h6 == idxUpdate_4[3:0]) begin
            TBEValid_6 <= 1'h0;
          end else begin
            TBEValid_6 <= _GEN_2045;
          end
        end else begin
          TBEValid_6 <= _GEN_2045;
        end
      end else if (isAlloc_4) begin
        TBEValid_6 <= _GEN_2126;
      end else if (_T_177) begin
        if (4'h6 == idxUpdate_4[3:0]) begin
          TBEValid_6 <= 1'h0;
        end else begin
          TBEValid_6 <= _GEN_2045;
        end
      end else begin
        TBEValid_6 <= _GEN_2045;
      end
    end else if (isAlloc_6) begin
      TBEValid_6 <= _GEN_3154;
    end else if (_T_221) begin
      if (4'h6 == idxUpdate_6[3:0]) begin
        TBEValid_6 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_6 <= _GEN_2640;
      end else if (_T_199) begin
        if (4'h6 == idxUpdate_5[3:0]) begin
          TBEValid_6 <= 1'h0;
        end else begin
          TBEValid_6 <= _GEN_2559;
        end
      end else begin
        TBEValid_6 <= _GEN_2559;
      end
    end else if (isAlloc_5) begin
      TBEValid_6 <= _GEN_2640;
    end else if (_T_199) begin
      if (4'h6 == idxUpdate_5[3:0]) begin
        TBEValid_6 <= 1'h0;
      end else begin
        TBEValid_6 <= _GEN_2559;
      end
    end else begin
      TBEValid_6 <= _GEN_2559;
    end
    if (reset) begin
      TBEValid_7 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_7 <= _GEN_3669;
    end else if (_T_243) begin
      if (4'h7 == idxUpdate_7[3:0]) begin
        TBEValid_7 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_7 <= _GEN_3155;
      end else if (_T_221) begin
        if (4'h7 == idxUpdate_6[3:0]) begin
          TBEValid_7 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_7 <= _GEN_2641;
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEValid_7 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_7 <= _GEN_2127;
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEValid_7 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_7 <= _GEN_1613;
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEValid_7 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_7 <= _GEN_1099;
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEValid_7 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_7 <= _GEN_585;
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEValid_7 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_7 <= _GEN_71;
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEValid_7 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_7 <= _GEN_71;
                end else if (_T_89) begin
                  if (4'h7 == idxUpdate_0[3:0]) begin
                    TBEValid_7 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_7 <= _GEN_585;
              end else if (_T_111) begin
                if (4'h7 == idxUpdate_1[3:0]) begin
                  TBEValid_7 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_7 <= _GEN_71;
                end else if (_T_89) begin
                  if (4'h7 == idxUpdate_0[3:0]) begin
                    TBEValid_7 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_7 <= _GEN_71;
              end else if (_T_89) begin
                if (4'h7 == idxUpdate_0[3:0]) begin
                  TBEValid_7 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_7 <= _GEN_1099;
            end else if (_T_133) begin
              if (4'h7 == idxUpdate_2[3:0]) begin
                TBEValid_7 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_7 <= _GEN_585;
              end else if (_T_111) begin
                if (4'h7 == idxUpdate_1[3:0]) begin
                  TBEValid_7 <= 1'h0;
                end else begin
                  TBEValid_7 <= _GEN_504;
                end
              end else begin
                TBEValid_7 <= _GEN_504;
              end
            end else if (isAlloc_1) begin
              TBEValid_7 <= _GEN_585;
            end else if (_T_111) begin
              if (4'h7 == idxUpdate_1[3:0]) begin
                TBEValid_7 <= 1'h0;
              end else begin
                TBEValid_7 <= _GEN_504;
              end
            end else begin
              TBEValid_7 <= _GEN_504;
            end
          end else if (isAlloc_3) begin
            TBEValid_7 <= _GEN_1613;
          end else if (_T_155) begin
            if (4'h7 == idxUpdate_3[3:0]) begin
              TBEValid_7 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_7 <= _GEN_1099;
            end else if (_T_133) begin
              if (4'h7 == idxUpdate_2[3:0]) begin
                TBEValid_7 <= 1'h0;
              end else begin
                TBEValid_7 <= _GEN_1018;
              end
            end else begin
              TBEValid_7 <= _GEN_1018;
            end
          end else if (isAlloc_2) begin
            TBEValid_7 <= _GEN_1099;
          end else if (_T_133) begin
            if (4'h7 == idxUpdate_2[3:0]) begin
              TBEValid_7 <= 1'h0;
            end else begin
              TBEValid_7 <= _GEN_1018;
            end
          end else begin
            TBEValid_7 <= _GEN_1018;
          end
        end else if (isAlloc_4) begin
          TBEValid_7 <= _GEN_2127;
        end else if (_T_177) begin
          if (4'h7 == idxUpdate_4[3:0]) begin
            TBEValid_7 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_7 <= _GEN_1613;
          end else if (_T_155) begin
            if (4'h7 == idxUpdate_3[3:0]) begin
              TBEValid_7 <= 1'h0;
            end else begin
              TBEValid_7 <= _GEN_1532;
            end
          end else begin
            TBEValid_7 <= _GEN_1532;
          end
        end else if (isAlloc_3) begin
          TBEValid_7 <= _GEN_1613;
        end else if (_T_155) begin
          if (4'h7 == idxUpdate_3[3:0]) begin
            TBEValid_7 <= 1'h0;
          end else begin
            TBEValid_7 <= _GEN_1532;
          end
        end else begin
          TBEValid_7 <= _GEN_1532;
        end
      end else if (isAlloc_5) begin
        TBEValid_7 <= _GEN_2641;
      end else if (_T_199) begin
        if (4'h7 == idxUpdate_5[3:0]) begin
          TBEValid_7 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_7 <= _GEN_2127;
        end else if (_T_177) begin
          if (4'h7 == idxUpdate_4[3:0]) begin
            TBEValid_7 <= 1'h0;
          end else begin
            TBEValid_7 <= _GEN_2046;
          end
        end else begin
          TBEValid_7 <= _GEN_2046;
        end
      end else if (isAlloc_4) begin
        TBEValid_7 <= _GEN_2127;
      end else if (_T_177) begin
        if (4'h7 == idxUpdate_4[3:0]) begin
          TBEValid_7 <= 1'h0;
        end else begin
          TBEValid_7 <= _GEN_2046;
        end
      end else begin
        TBEValid_7 <= _GEN_2046;
      end
    end else if (isAlloc_6) begin
      TBEValid_7 <= _GEN_3155;
    end else if (_T_221) begin
      if (4'h7 == idxUpdate_6[3:0]) begin
        TBEValid_7 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_7 <= _GEN_2641;
      end else if (_T_199) begin
        if (4'h7 == idxUpdate_5[3:0]) begin
          TBEValid_7 <= 1'h0;
        end else begin
          TBEValid_7 <= _GEN_2560;
        end
      end else begin
        TBEValid_7 <= _GEN_2560;
      end
    end else if (isAlloc_5) begin
      TBEValid_7 <= _GEN_2641;
    end else if (_T_199) begin
      if (4'h7 == idxUpdate_5[3:0]) begin
        TBEValid_7 <= 1'h0;
      end else begin
        TBEValid_7 <= _GEN_2560;
      end
    end else begin
      TBEValid_7 <= _GEN_2560;
    end
    if (reset) begin
      TBEValid_8 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_8 <= _GEN_3670;
    end else if (_T_243) begin
      if (4'h8 == idxUpdate_7[3:0]) begin
        TBEValid_8 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_8 <= _GEN_3156;
      end else if (_T_221) begin
        if (4'h8 == idxUpdate_6[3:0]) begin
          TBEValid_8 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_8 <= _GEN_2642;
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEValid_8 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_8 <= _GEN_2128;
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEValid_8 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_8 <= _GEN_1614;
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEValid_8 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_8 <= _GEN_1100;
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEValid_8 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_8 <= _GEN_586;
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEValid_8 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_8 <= _GEN_72;
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEValid_8 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_8 <= _GEN_72;
                end else if (_T_89) begin
                  if (4'h8 == idxUpdate_0[3:0]) begin
                    TBEValid_8 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_8 <= _GEN_586;
              end else if (_T_111) begin
                if (4'h8 == idxUpdate_1[3:0]) begin
                  TBEValid_8 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_8 <= _GEN_72;
                end else if (_T_89) begin
                  if (4'h8 == idxUpdate_0[3:0]) begin
                    TBEValid_8 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_8 <= _GEN_72;
              end else if (_T_89) begin
                if (4'h8 == idxUpdate_0[3:0]) begin
                  TBEValid_8 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_8 <= _GEN_1100;
            end else if (_T_133) begin
              if (4'h8 == idxUpdate_2[3:0]) begin
                TBEValid_8 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_8 <= _GEN_586;
              end else if (_T_111) begin
                if (4'h8 == idxUpdate_1[3:0]) begin
                  TBEValid_8 <= 1'h0;
                end else begin
                  TBEValid_8 <= _GEN_505;
                end
              end else begin
                TBEValid_8 <= _GEN_505;
              end
            end else if (isAlloc_1) begin
              TBEValid_8 <= _GEN_586;
            end else if (_T_111) begin
              if (4'h8 == idxUpdate_1[3:0]) begin
                TBEValid_8 <= 1'h0;
              end else begin
                TBEValid_8 <= _GEN_505;
              end
            end else begin
              TBEValid_8 <= _GEN_505;
            end
          end else if (isAlloc_3) begin
            TBEValid_8 <= _GEN_1614;
          end else if (_T_155) begin
            if (4'h8 == idxUpdate_3[3:0]) begin
              TBEValid_8 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_8 <= _GEN_1100;
            end else if (_T_133) begin
              if (4'h8 == idxUpdate_2[3:0]) begin
                TBEValid_8 <= 1'h0;
              end else begin
                TBEValid_8 <= _GEN_1019;
              end
            end else begin
              TBEValid_8 <= _GEN_1019;
            end
          end else if (isAlloc_2) begin
            TBEValid_8 <= _GEN_1100;
          end else if (_T_133) begin
            if (4'h8 == idxUpdate_2[3:0]) begin
              TBEValid_8 <= 1'h0;
            end else begin
              TBEValid_8 <= _GEN_1019;
            end
          end else begin
            TBEValid_8 <= _GEN_1019;
          end
        end else if (isAlloc_4) begin
          TBEValid_8 <= _GEN_2128;
        end else if (_T_177) begin
          if (4'h8 == idxUpdate_4[3:0]) begin
            TBEValid_8 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_8 <= _GEN_1614;
          end else if (_T_155) begin
            if (4'h8 == idxUpdate_3[3:0]) begin
              TBEValid_8 <= 1'h0;
            end else begin
              TBEValid_8 <= _GEN_1533;
            end
          end else begin
            TBEValid_8 <= _GEN_1533;
          end
        end else if (isAlloc_3) begin
          TBEValid_8 <= _GEN_1614;
        end else if (_T_155) begin
          if (4'h8 == idxUpdate_3[3:0]) begin
            TBEValid_8 <= 1'h0;
          end else begin
            TBEValid_8 <= _GEN_1533;
          end
        end else begin
          TBEValid_8 <= _GEN_1533;
        end
      end else if (isAlloc_5) begin
        TBEValid_8 <= _GEN_2642;
      end else if (_T_199) begin
        if (4'h8 == idxUpdate_5[3:0]) begin
          TBEValid_8 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_8 <= _GEN_2128;
        end else if (_T_177) begin
          if (4'h8 == idxUpdate_4[3:0]) begin
            TBEValid_8 <= 1'h0;
          end else begin
            TBEValid_8 <= _GEN_2047;
          end
        end else begin
          TBEValid_8 <= _GEN_2047;
        end
      end else if (isAlloc_4) begin
        TBEValid_8 <= _GEN_2128;
      end else if (_T_177) begin
        if (4'h8 == idxUpdate_4[3:0]) begin
          TBEValid_8 <= 1'h0;
        end else begin
          TBEValid_8 <= _GEN_2047;
        end
      end else begin
        TBEValid_8 <= _GEN_2047;
      end
    end else if (isAlloc_6) begin
      TBEValid_8 <= _GEN_3156;
    end else if (_T_221) begin
      if (4'h8 == idxUpdate_6[3:0]) begin
        TBEValid_8 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_8 <= _GEN_2642;
      end else if (_T_199) begin
        if (4'h8 == idxUpdate_5[3:0]) begin
          TBEValid_8 <= 1'h0;
        end else begin
          TBEValid_8 <= _GEN_2561;
        end
      end else begin
        TBEValid_8 <= _GEN_2561;
      end
    end else if (isAlloc_5) begin
      TBEValid_8 <= _GEN_2642;
    end else if (_T_199) begin
      if (4'h8 == idxUpdate_5[3:0]) begin
        TBEValid_8 <= 1'h0;
      end else begin
        TBEValid_8 <= _GEN_2561;
      end
    end else begin
      TBEValid_8 <= _GEN_2561;
    end
    if (reset) begin
      TBEValid_9 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_9 <= _GEN_3671;
    end else if (_T_243) begin
      if (4'h9 == idxUpdate_7[3:0]) begin
        TBEValid_9 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_9 <= _GEN_3157;
      end else if (_T_221) begin
        if (4'h9 == idxUpdate_6[3:0]) begin
          TBEValid_9 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_9 <= _GEN_2643;
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEValid_9 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_9 <= _GEN_2129;
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEValid_9 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_9 <= _GEN_1615;
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEValid_9 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_9 <= _GEN_1101;
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEValid_9 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_9 <= _GEN_587;
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEValid_9 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_9 <= _GEN_73;
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEValid_9 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_9 <= _GEN_73;
                end else if (_T_89) begin
                  if (4'h9 == idxUpdate_0[3:0]) begin
                    TBEValid_9 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_9 <= _GEN_587;
              end else if (_T_111) begin
                if (4'h9 == idxUpdate_1[3:0]) begin
                  TBEValid_9 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_9 <= _GEN_73;
                end else if (_T_89) begin
                  if (4'h9 == idxUpdate_0[3:0]) begin
                    TBEValid_9 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_9 <= _GEN_73;
              end else if (_T_89) begin
                if (4'h9 == idxUpdate_0[3:0]) begin
                  TBEValid_9 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_9 <= _GEN_1101;
            end else if (_T_133) begin
              if (4'h9 == idxUpdate_2[3:0]) begin
                TBEValid_9 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_9 <= _GEN_587;
              end else if (_T_111) begin
                if (4'h9 == idxUpdate_1[3:0]) begin
                  TBEValid_9 <= 1'h0;
                end else begin
                  TBEValid_9 <= _GEN_506;
                end
              end else begin
                TBEValid_9 <= _GEN_506;
              end
            end else if (isAlloc_1) begin
              TBEValid_9 <= _GEN_587;
            end else if (_T_111) begin
              if (4'h9 == idxUpdate_1[3:0]) begin
                TBEValid_9 <= 1'h0;
              end else begin
                TBEValid_9 <= _GEN_506;
              end
            end else begin
              TBEValid_9 <= _GEN_506;
            end
          end else if (isAlloc_3) begin
            TBEValid_9 <= _GEN_1615;
          end else if (_T_155) begin
            if (4'h9 == idxUpdate_3[3:0]) begin
              TBEValid_9 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_9 <= _GEN_1101;
            end else if (_T_133) begin
              if (4'h9 == idxUpdate_2[3:0]) begin
                TBEValid_9 <= 1'h0;
              end else begin
                TBEValid_9 <= _GEN_1020;
              end
            end else begin
              TBEValid_9 <= _GEN_1020;
            end
          end else if (isAlloc_2) begin
            TBEValid_9 <= _GEN_1101;
          end else if (_T_133) begin
            if (4'h9 == idxUpdate_2[3:0]) begin
              TBEValid_9 <= 1'h0;
            end else begin
              TBEValid_9 <= _GEN_1020;
            end
          end else begin
            TBEValid_9 <= _GEN_1020;
          end
        end else if (isAlloc_4) begin
          TBEValid_9 <= _GEN_2129;
        end else if (_T_177) begin
          if (4'h9 == idxUpdate_4[3:0]) begin
            TBEValid_9 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_9 <= _GEN_1615;
          end else if (_T_155) begin
            if (4'h9 == idxUpdate_3[3:0]) begin
              TBEValid_9 <= 1'h0;
            end else begin
              TBEValid_9 <= _GEN_1534;
            end
          end else begin
            TBEValid_9 <= _GEN_1534;
          end
        end else if (isAlloc_3) begin
          TBEValid_9 <= _GEN_1615;
        end else if (_T_155) begin
          if (4'h9 == idxUpdate_3[3:0]) begin
            TBEValid_9 <= 1'h0;
          end else begin
            TBEValid_9 <= _GEN_1534;
          end
        end else begin
          TBEValid_9 <= _GEN_1534;
        end
      end else if (isAlloc_5) begin
        TBEValid_9 <= _GEN_2643;
      end else if (_T_199) begin
        if (4'h9 == idxUpdate_5[3:0]) begin
          TBEValid_9 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_9 <= _GEN_2129;
        end else if (_T_177) begin
          if (4'h9 == idxUpdate_4[3:0]) begin
            TBEValid_9 <= 1'h0;
          end else begin
            TBEValid_9 <= _GEN_2048;
          end
        end else begin
          TBEValid_9 <= _GEN_2048;
        end
      end else if (isAlloc_4) begin
        TBEValid_9 <= _GEN_2129;
      end else if (_T_177) begin
        if (4'h9 == idxUpdate_4[3:0]) begin
          TBEValid_9 <= 1'h0;
        end else begin
          TBEValid_9 <= _GEN_2048;
        end
      end else begin
        TBEValid_9 <= _GEN_2048;
      end
    end else if (isAlloc_6) begin
      TBEValid_9 <= _GEN_3157;
    end else if (_T_221) begin
      if (4'h9 == idxUpdate_6[3:0]) begin
        TBEValid_9 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_9 <= _GEN_2643;
      end else if (_T_199) begin
        if (4'h9 == idxUpdate_5[3:0]) begin
          TBEValid_9 <= 1'h0;
        end else begin
          TBEValid_9 <= _GEN_2562;
        end
      end else begin
        TBEValid_9 <= _GEN_2562;
      end
    end else if (isAlloc_5) begin
      TBEValid_9 <= _GEN_2643;
    end else if (_T_199) begin
      if (4'h9 == idxUpdate_5[3:0]) begin
        TBEValid_9 <= 1'h0;
      end else begin
        TBEValid_9 <= _GEN_2562;
      end
    end else begin
      TBEValid_9 <= _GEN_2562;
    end
    if (reset) begin
      TBEValid_10 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_10 <= _GEN_3672;
    end else if (_T_243) begin
      if (4'ha == idxUpdate_7[3:0]) begin
        TBEValid_10 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_10 <= _GEN_3158;
      end else if (_T_221) begin
        if (4'ha == idxUpdate_6[3:0]) begin
          TBEValid_10 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_10 <= _GEN_2644;
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEValid_10 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_10 <= _GEN_2130;
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEValid_10 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_10 <= _GEN_1616;
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEValid_10 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_10 <= _GEN_1102;
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEValid_10 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_10 <= _GEN_588;
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEValid_10 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_10 <= _GEN_74;
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEValid_10 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_10 <= _GEN_74;
                end else if (_T_89) begin
                  if (4'ha == idxUpdate_0[3:0]) begin
                    TBEValid_10 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_10 <= _GEN_588;
              end else if (_T_111) begin
                if (4'ha == idxUpdate_1[3:0]) begin
                  TBEValid_10 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_10 <= _GEN_74;
                end else if (_T_89) begin
                  if (4'ha == idxUpdate_0[3:0]) begin
                    TBEValid_10 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_10 <= _GEN_74;
              end else if (_T_89) begin
                if (4'ha == idxUpdate_0[3:0]) begin
                  TBEValid_10 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_10 <= _GEN_1102;
            end else if (_T_133) begin
              if (4'ha == idxUpdate_2[3:0]) begin
                TBEValid_10 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_10 <= _GEN_588;
              end else if (_T_111) begin
                if (4'ha == idxUpdate_1[3:0]) begin
                  TBEValid_10 <= 1'h0;
                end else begin
                  TBEValid_10 <= _GEN_507;
                end
              end else begin
                TBEValid_10 <= _GEN_507;
              end
            end else if (isAlloc_1) begin
              TBEValid_10 <= _GEN_588;
            end else if (_T_111) begin
              if (4'ha == idxUpdate_1[3:0]) begin
                TBEValid_10 <= 1'h0;
              end else begin
                TBEValid_10 <= _GEN_507;
              end
            end else begin
              TBEValid_10 <= _GEN_507;
            end
          end else if (isAlloc_3) begin
            TBEValid_10 <= _GEN_1616;
          end else if (_T_155) begin
            if (4'ha == idxUpdate_3[3:0]) begin
              TBEValid_10 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_10 <= _GEN_1102;
            end else if (_T_133) begin
              if (4'ha == idxUpdate_2[3:0]) begin
                TBEValid_10 <= 1'h0;
              end else begin
                TBEValid_10 <= _GEN_1021;
              end
            end else begin
              TBEValid_10 <= _GEN_1021;
            end
          end else if (isAlloc_2) begin
            TBEValid_10 <= _GEN_1102;
          end else if (_T_133) begin
            if (4'ha == idxUpdate_2[3:0]) begin
              TBEValid_10 <= 1'h0;
            end else begin
              TBEValid_10 <= _GEN_1021;
            end
          end else begin
            TBEValid_10 <= _GEN_1021;
          end
        end else if (isAlloc_4) begin
          TBEValid_10 <= _GEN_2130;
        end else if (_T_177) begin
          if (4'ha == idxUpdate_4[3:0]) begin
            TBEValid_10 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_10 <= _GEN_1616;
          end else if (_T_155) begin
            if (4'ha == idxUpdate_3[3:0]) begin
              TBEValid_10 <= 1'h0;
            end else begin
              TBEValid_10 <= _GEN_1535;
            end
          end else begin
            TBEValid_10 <= _GEN_1535;
          end
        end else if (isAlloc_3) begin
          TBEValid_10 <= _GEN_1616;
        end else if (_T_155) begin
          if (4'ha == idxUpdate_3[3:0]) begin
            TBEValid_10 <= 1'h0;
          end else begin
            TBEValid_10 <= _GEN_1535;
          end
        end else begin
          TBEValid_10 <= _GEN_1535;
        end
      end else if (isAlloc_5) begin
        TBEValid_10 <= _GEN_2644;
      end else if (_T_199) begin
        if (4'ha == idxUpdate_5[3:0]) begin
          TBEValid_10 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_10 <= _GEN_2130;
        end else if (_T_177) begin
          if (4'ha == idxUpdate_4[3:0]) begin
            TBEValid_10 <= 1'h0;
          end else begin
            TBEValid_10 <= _GEN_2049;
          end
        end else begin
          TBEValid_10 <= _GEN_2049;
        end
      end else if (isAlloc_4) begin
        TBEValid_10 <= _GEN_2130;
      end else if (_T_177) begin
        if (4'ha == idxUpdate_4[3:0]) begin
          TBEValid_10 <= 1'h0;
        end else begin
          TBEValid_10 <= _GEN_2049;
        end
      end else begin
        TBEValid_10 <= _GEN_2049;
      end
    end else if (isAlloc_6) begin
      TBEValid_10 <= _GEN_3158;
    end else if (_T_221) begin
      if (4'ha == idxUpdate_6[3:0]) begin
        TBEValid_10 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_10 <= _GEN_2644;
      end else if (_T_199) begin
        if (4'ha == idxUpdate_5[3:0]) begin
          TBEValid_10 <= 1'h0;
        end else begin
          TBEValid_10 <= _GEN_2563;
        end
      end else begin
        TBEValid_10 <= _GEN_2563;
      end
    end else if (isAlloc_5) begin
      TBEValid_10 <= _GEN_2644;
    end else if (_T_199) begin
      if (4'ha == idxUpdate_5[3:0]) begin
        TBEValid_10 <= 1'h0;
      end else begin
        TBEValid_10 <= _GEN_2563;
      end
    end else begin
      TBEValid_10 <= _GEN_2563;
    end
    if (reset) begin
      TBEValid_11 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_11 <= _GEN_3673;
    end else if (_T_243) begin
      if (4'hb == idxUpdate_7[3:0]) begin
        TBEValid_11 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_11 <= _GEN_3159;
      end else if (_T_221) begin
        if (4'hb == idxUpdate_6[3:0]) begin
          TBEValid_11 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_11 <= _GEN_2645;
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEValid_11 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_11 <= _GEN_2131;
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEValid_11 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_11 <= _GEN_1617;
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEValid_11 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_11 <= _GEN_1103;
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEValid_11 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_11 <= _GEN_589;
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEValid_11 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_11 <= _GEN_75;
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEValid_11 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_11 <= _GEN_75;
                end else if (_T_89) begin
                  if (4'hb == idxUpdate_0[3:0]) begin
                    TBEValid_11 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_11 <= _GEN_589;
              end else if (_T_111) begin
                if (4'hb == idxUpdate_1[3:0]) begin
                  TBEValid_11 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_11 <= _GEN_75;
                end else if (_T_89) begin
                  if (4'hb == idxUpdate_0[3:0]) begin
                    TBEValid_11 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_11 <= _GEN_75;
              end else if (_T_89) begin
                if (4'hb == idxUpdate_0[3:0]) begin
                  TBEValid_11 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_11 <= _GEN_1103;
            end else if (_T_133) begin
              if (4'hb == idxUpdate_2[3:0]) begin
                TBEValid_11 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_11 <= _GEN_589;
              end else if (_T_111) begin
                if (4'hb == idxUpdate_1[3:0]) begin
                  TBEValid_11 <= 1'h0;
                end else begin
                  TBEValid_11 <= _GEN_508;
                end
              end else begin
                TBEValid_11 <= _GEN_508;
              end
            end else if (isAlloc_1) begin
              TBEValid_11 <= _GEN_589;
            end else if (_T_111) begin
              if (4'hb == idxUpdate_1[3:0]) begin
                TBEValid_11 <= 1'h0;
              end else begin
                TBEValid_11 <= _GEN_508;
              end
            end else begin
              TBEValid_11 <= _GEN_508;
            end
          end else if (isAlloc_3) begin
            TBEValid_11 <= _GEN_1617;
          end else if (_T_155) begin
            if (4'hb == idxUpdate_3[3:0]) begin
              TBEValid_11 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_11 <= _GEN_1103;
            end else if (_T_133) begin
              if (4'hb == idxUpdate_2[3:0]) begin
                TBEValid_11 <= 1'h0;
              end else begin
                TBEValid_11 <= _GEN_1022;
              end
            end else begin
              TBEValid_11 <= _GEN_1022;
            end
          end else if (isAlloc_2) begin
            TBEValid_11 <= _GEN_1103;
          end else if (_T_133) begin
            if (4'hb == idxUpdate_2[3:0]) begin
              TBEValid_11 <= 1'h0;
            end else begin
              TBEValid_11 <= _GEN_1022;
            end
          end else begin
            TBEValid_11 <= _GEN_1022;
          end
        end else if (isAlloc_4) begin
          TBEValid_11 <= _GEN_2131;
        end else if (_T_177) begin
          if (4'hb == idxUpdate_4[3:0]) begin
            TBEValid_11 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_11 <= _GEN_1617;
          end else if (_T_155) begin
            if (4'hb == idxUpdate_3[3:0]) begin
              TBEValid_11 <= 1'h0;
            end else begin
              TBEValid_11 <= _GEN_1536;
            end
          end else begin
            TBEValid_11 <= _GEN_1536;
          end
        end else if (isAlloc_3) begin
          TBEValid_11 <= _GEN_1617;
        end else if (_T_155) begin
          if (4'hb == idxUpdate_3[3:0]) begin
            TBEValid_11 <= 1'h0;
          end else begin
            TBEValid_11 <= _GEN_1536;
          end
        end else begin
          TBEValid_11 <= _GEN_1536;
        end
      end else if (isAlloc_5) begin
        TBEValid_11 <= _GEN_2645;
      end else if (_T_199) begin
        if (4'hb == idxUpdate_5[3:0]) begin
          TBEValid_11 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_11 <= _GEN_2131;
        end else if (_T_177) begin
          if (4'hb == idxUpdate_4[3:0]) begin
            TBEValid_11 <= 1'h0;
          end else begin
            TBEValid_11 <= _GEN_2050;
          end
        end else begin
          TBEValid_11 <= _GEN_2050;
        end
      end else if (isAlloc_4) begin
        TBEValid_11 <= _GEN_2131;
      end else if (_T_177) begin
        if (4'hb == idxUpdate_4[3:0]) begin
          TBEValid_11 <= 1'h0;
        end else begin
          TBEValid_11 <= _GEN_2050;
        end
      end else begin
        TBEValid_11 <= _GEN_2050;
      end
    end else if (isAlloc_6) begin
      TBEValid_11 <= _GEN_3159;
    end else if (_T_221) begin
      if (4'hb == idxUpdate_6[3:0]) begin
        TBEValid_11 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_11 <= _GEN_2645;
      end else if (_T_199) begin
        if (4'hb == idxUpdate_5[3:0]) begin
          TBEValid_11 <= 1'h0;
        end else begin
          TBEValid_11 <= _GEN_2564;
        end
      end else begin
        TBEValid_11 <= _GEN_2564;
      end
    end else if (isAlloc_5) begin
      TBEValid_11 <= _GEN_2645;
    end else if (_T_199) begin
      if (4'hb == idxUpdate_5[3:0]) begin
        TBEValid_11 <= 1'h0;
      end else begin
        TBEValid_11 <= _GEN_2564;
      end
    end else begin
      TBEValid_11 <= _GEN_2564;
    end
    if (reset) begin
      TBEValid_12 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_12 <= _GEN_3674;
    end else if (_T_243) begin
      if (4'hc == idxUpdate_7[3:0]) begin
        TBEValid_12 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_12 <= _GEN_3160;
      end else if (_T_221) begin
        if (4'hc == idxUpdate_6[3:0]) begin
          TBEValid_12 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_12 <= _GEN_2646;
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEValid_12 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_12 <= _GEN_2132;
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEValid_12 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_12 <= _GEN_1618;
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEValid_12 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_12 <= _GEN_1104;
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEValid_12 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_12 <= _GEN_590;
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEValid_12 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_12 <= _GEN_76;
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEValid_12 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_12 <= _GEN_76;
                end else if (_T_89) begin
                  if (4'hc == idxUpdate_0[3:0]) begin
                    TBEValid_12 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_12 <= _GEN_590;
              end else if (_T_111) begin
                if (4'hc == idxUpdate_1[3:0]) begin
                  TBEValid_12 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_12 <= _GEN_76;
                end else if (_T_89) begin
                  if (4'hc == idxUpdate_0[3:0]) begin
                    TBEValid_12 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_12 <= _GEN_76;
              end else if (_T_89) begin
                if (4'hc == idxUpdate_0[3:0]) begin
                  TBEValid_12 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_12 <= _GEN_1104;
            end else if (_T_133) begin
              if (4'hc == idxUpdate_2[3:0]) begin
                TBEValid_12 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_12 <= _GEN_590;
              end else if (_T_111) begin
                if (4'hc == idxUpdate_1[3:0]) begin
                  TBEValid_12 <= 1'h0;
                end else begin
                  TBEValid_12 <= _GEN_509;
                end
              end else begin
                TBEValid_12 <= _GEN_509;
              end
            end else if (isAlloc_1) begin
              TBEValid_12 <= _GEN_590;
            end else if (_T_111) begin
              if (4'hc == idxUpdate_1[3:0]) begin
                TBEValid_12 <= 1'h0;
              end else begin
                TBEValid_12 <= _GEN_509;
              end
            end else begin
              TBEValid_12 <= _GEN_509;
            end
          end else if (isAlloc_3) begin
            TBEValid_12 <= _GEN_1618;
          end else if (_T_155) begin
            if (4'hc == idxUpdate_3[3:0]) begin
              TBEValid_12 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_12 <= _GEN_1104;
            end else if (_T_133) begin
              if (4'hc == idxUpdate_2[3:0]) begin
                TBEValid_12 <= 1'h0;
              end else begin
                TBEValid_12 <= _GEN_1023;
              end
            end else begin
              TBEValid_12 <= _GEN_1023;
            end
          end else if (isAlloc_2) begin
            TBEValid_12 <= _GEN_1104;
          end else if (_T_133) begin
            if (4'hc == idxUpdate_2[3:0]) begin
              TBEValid_12 <= 1'h0;
            end else begin
              TBEValid_12 <= _GEN_1023;
            end
          end else begin
            TBEValid_12 <= _GEN_1023;
          end
        end else if (isAlloc_4) begin
          TBEValid_12 <= _GEN_2132;
        end else if (_T_177) begin
          if (4'hc == idxUpdate_4[3:0]) begin
            TBEValid_12 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_12 <= _GEN_1618;
          end else if (_T_155) begin
            if (4'hc == idxUpdate_3[3:0]) begin
              TBEValid_12 <= 1'h0;
            end else begin
              TBEValid_12 <= _GEN_1537;
            end
          end else begin
            TBEValid_12 <= _GEN_1537;
          end
        end else if (isAlloc_3) begin
          TBEValid_12 <= _GEN_1618;
        end else if (_T_155) begin
          if (4'hc == idxUpdate_3[3:0]) begin
            TBEValid_12 <= 1'h0;
          end else begin
            TBEValid_12 <= _GEN_1537;
          end
        end else begin
          TBEValid_12 <= _GEN_1537;
        end
      end else if (isAlloc_5) begin
        TBEValid_12 <= _GEN_2646;
      end else if (_T_199) begin
        if (4'hc == idxUpdate_5[3:0]) begin
          TBEValid_12 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_12 <= _GEN_2132;
        end else if (_T_177) begin
          if (4'hc == idxUpdate_4[3:0]) begin
            TBEValid_12 <= 1'h0;
          end else begin
            TBEValid_12 <= _GEN_2051;
          end
        end else begin
          TBEValid_12 <= _GEN_2051;
        end
      end else if (isAlloc_4) begin
        TBEValid_12 <= _GEN_2132;
      end else if (_T_177) begin
        if (4'hc == idxUpdate_4[3:0]) begin
          TBEValid_12 <= 1'h0;
        end else begin
          TBEValid_12 <= _GEN_2051;
        end
      end else begin
        TBEValid_12 <= _GEN_2051;
      end
    end else if (isAlloc_6) begin
      TBEValid_12 <= _GEN_3160;
    end else if (_T_221) begin
      if (4'hc == idxUpdate_6[3:0]) begin
        TBEValid_12 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_12 <= _GEN_2646;
      end else if (_T_199) begin
        if (4'hc == idxUpdate_5[3:0]) begin
          TBEValid_12 <= 1'h0;
        end else begin
          TBEValid_12 <= _GEN_2565;
        end
      end else begin
        TBEValid_12 <= _GEN_2565;
      end
    end else if (isAlloc_5) begin
      TBEValid_12 <= _GEN_2646;
    end else if (_T_199) begin
      if (4'hc == idxUpdate_5[3:0]) begin
        TBEValid_12 <= 1'h0;
      end else begin
        TBEValid_12 <= _GEN_2565;
      end
    end else begin
      TBEValid_12 <= _GEN_2565;
    end
    if (reset) begin
      TBEValid_13 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_13 <= _GEN_3675;
    end else if (_T_243) begin
      if (4'hd == idxUpdate_7[3:0]) begin
        TBEValid_13 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_13 <= _GEN_3161;
      end else if (_T_221) begin
        if (4'hd == idxUpdate_6[3:0]) begin
          TBEValid_13 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_13 <= _GEN_2647;
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEValid_13 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_13 <= _GEN_2133;
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEValid_13 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_13 <= _GEN_1619;
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEValid_13 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_13 <= _GEN_1105;
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEValid_13 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_13 <= _GEN_591;
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEValid_13 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_13 <= _GEN_77;
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEValid_13 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_13 <= _GEN_77;
                end else if (_T_89) begin
                  if (4'hd == idxUpdate_0[3:0]) begin
                    TBEValid_13 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_13 <= _GEN_591;
              end else if (_T_111) begin
                if (4'hd == idxUpdate_1[3:0]) begin
                  TBEValid_13 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_13 <= _GEN_77;
                end else if (_T_89) begin
                  if (4'hd == idxUpdate_0[3:0]) begin
                    TBEValid_13 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_13 <= _GEN_77;
              end else if (_T_89) begin
                if (4'hd == idxUpdate_0[3:0]) begin
                  TBEValid_13 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_13 <= _GEN_1105;
            end else if (_T_133) begin
              if (4'hd == idxUpdate_2[3:0]) begin
                TBEValid_13 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_13 <= _GEN_591;
              end else if (_T_111) begin
                if (4'hd == idxUpdate_1[3:0]) begin
                  TBEValid_13 <= 1'h0;
                end else begin
                  TBEValid_13 <= _GEN_510;
                end
              end else begin
                TBEValid_13 <= _GEN_510;
              end
            end else if (isAlloc_1) begin
              TBEValid_13 <= _GEN_591;
            end else if (_T_111) begin
              if (4'hd == idxUpdate_1[3:0]) begin
                TBEValid_13 <= 1'h0;
              end else begin
                TBEValid_13 <= _GEN_510;
              end
            end else begin
              TBEValid_13 <= _GEN_510;
            end
          end else if (isAlloc_3) begin
            TBEValid_13 <= _GEN_1619;
          end else if (_T_155) begin
            if (4'hd == idxUpdate_3[3:0]) begin
              TBEValid_13 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_13 <= _GEN_1105;
            end else if (_T_133) begin
              if (4'hd == idxUpdate_2[3:0]) begin
                TBEValid_13 <= 1'h0;
              end else begin
                TBEValid_13 <= _GEN_1024;
              end
            end else begin
              TBEValid_13 <= _GEN_1024;
            end
          end else if (isAlloc_2) begin
            TBEValid_13 <= _GEN_1105;
          end else if (_T_133) begin
            if (4'hd == idxUpdate_2[3:0]) begin
              TBEValid_13 <= 1'h0;
            end else begin
              TBEValid_13 <= _GEN_1024;
            end
          end else begin
            TBEValid_13 <= _GEN_1024;
          end
        end else if (isAlloc_4) begin
          TBEValid_13 <= _GEN_2133;
        end else if (_T_177) begin
          if (4'hd == idxUpdate_4[3:0]) begin
            TBEValid_13 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_13 <= _GEN_1619;
          end else if (_T_155) begin
            if (4'hd == idxUpdate_3[3:0]) begin
              TBEValid_13 <= 1'h0;
            end else begin
              TBEValid_13 <= _GEN_1538;
            end
          end else begin
            TBEValid_13 <= _GEN_1538;
          end
        end else if (isAlloc_3) begin
          TBEValid_13 <= _GEN_1619;
        end else if (_T_155) begin
          if (4'hd == idxUpdate_3[3:0]) begin
            TBEValid_13 <= 1'h0;
          end else begin
            TBEValid_13 <= _GEN_1538;
          end
        end else begin
          TBEValid_13 <= _GEN_1538;
        end
      end else if (isAlloc_5) begin
        TBEValid_13 <= _GEN_2647;
      end else if (_T_199) begin
        if (4'hd == idxUpdate_5[3:0]) begin
          TBEValid_13 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_13 <= _GEN_2133;
        end else if (_T_177) begin
          if (4'hd == idxUpdate_4[3:0]) begin
            TBEValid_13 <= 1'h0;
          end else begin
            TBEValid_13 <= _GEN_2052;
          end
        end else begin
          TBEValid_13 <= _GEN_2052;
        end
      end else if (isAlloc_4) begin
        TBEValid_13 <= _GEN_2133;
      end else if (_T_177) begin
        if (4'hd == idxUpdate_4[3:0]) begin
          TBEValid_13 <= 1'h0;
        end else begin
          TBEValid_13 <= _GEN_2052;
        end
      end else begin
        TBEValid_13 <= _GEN_2052;
      end
    end else if (isAlloc_6) begin
      TBEValid_13 <= _GEN_3161;
    end else if (_T_221) begin
      if (4'hd == idxUpdate_6[3:0]) begin
        TBEValid_13 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_13 <= _GEN_2647;
      end else if (_T_199) begin
        if (4'hd == idxUpdate_5[3:0]) begin
          TBEValid_13 <= 1'h0;
        end else begin
          TBEValid_13 <= _GEN_2566;
        end
      end else begin
        TBEValid_13 <= _GEN_2566;
      end
    end else if (isAlloc_5) begin
      TBEValid_13 <= _GEN_2647;
    end else if (_T_199) begin
      if (4'hd == idxUpdate_5[3:0]) begin
        TBEValid_13 <= 1'h0;
      end else begin
        TBEValid_13 <= _GEN_2566;
      end
    end else begin
      TBEValid_13 <= _GEN_2566;
    end
    if (reset) begin
      TBEValid_14 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_14 <= _GEN_3676;
    end else if (_T_243) begin
      if (4'he == idxUpdate_7[3:0]) begin
        TBEValid_14 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_14 <= _GEN_3162;
      end else if (_T_221) begin
        if (4'he == idxUpdate_6[3:0]) begin
          TBEValid_14 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_14 <= _GEN_2648;
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEValid_14 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_14 <= _GEN_2134;
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEValid_14 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_14 <= _GEN_1620;
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEValid_14 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_14 <= _GEN_1106;
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEValid_14 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_14 <= _GEN_592;
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEValid_14 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_14 <= _GEN_78;
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEValid_14 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_14 <= _GEN_78;
                end else if (_T_89) begin
                  if (4'he == idxUpdate_0[3:0]) begin
                    TBEValid_14 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_14 <= _GEN_592;
              end else if (_T_111) begin
                if (4'he == idxUpdate_1[3:0]) begin
                  TBEValid_14 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_14 <= _GEN_78;
                end else if (_T_89) begin
                  if (4'he == idxUpdate_0[3:0]) begin
                    TBEValid_14 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_14 <= _GEN_78;
              end else if (_T_89) begin
                if (4'he == idxUpdate_0[3:0]) begin
                  TBEValid_14 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_14 <= _GEN_1106;
            end else if (_T_133) begin
              if (4'he == idxUpdate_2[3:0]) begin
                TBEValid_14 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_14 <= _GEN_592;
              end else if (_T_111) begin
                if (4'he == idxUpdate_1[3:0]) begin
                  TBEValid_14 <= 1'h0;
                end else begin
                  TBEValid_14 <= _GEN_511;
                end
              end else begin
                TBEValid_14 <= _GEN_511;
              end
            end else if (isAlloc_1) begin
              TBEValid_14 <= _GEN_592;
            end else if (_T_111) begin
              if (4'he == idxUpdate_1[3:0]) begin
                TBEValid_14 <= 1'h0;
              end else begin
                TBEValid_14 <= _GEN_511;
              end
            end else begin
              TBEValid_14 <= _GEN_511;
            end
          end else if (isAlloc_3) begin
            TBEValid_14 <= _GEN_1620;
          end else if (_T_155) begin
            if (4'he == idxUpdate_3[3:0]) begin
              TBEValid_14 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_14 <= _GEN_1106;
            end else if (_T_133) begin
              if (4'he == idxUpdate_2[3:0]) begin
                TBEValid_14 <= 1'h0;
              end else begin
                TBEValid_14 <= _GEN_1025;
              end
            end else begin
              TBEValid_14 <= _GEN_1025;
            end
          end else if (isAlloc_2) begin
            TBEValid_14 <= _GEN_1106;
          end else if (_T_133) begin
            if (4'he == idxUpdate_2[3:0]) begin
              TBEValid_14 <= 1'h0;
            end else begin
              TBEValid_14 <= _GEN_1025;
            end
          end else begin
            TBEValid_14 <= _GEN_1025;
          end
        end else if (isAlloc_4) begin
          TBEValid_14 <= _GEN_2134;
        end else if (_T_177) begin
          if (4'he == idxUpdate_4[3:0]) begin
            TBEValid_14 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_14 <= _GEN_1620;
          end else if (_T_155) begin
            if (4'he == idxUpdate_3[3:0]) begin
              TBEValid_14 <= 1'h0;
            end else begin
              TBEValid_14 <= _GEN_1539;
            end
          end else begin
            TBEValid_14 <= _GEN_1539;
          end
        end else if (isAlloc_3) begin
          TBEValid_14 <= _GEN_1620;
        end else if (_T_155) begin
          if (4'he == idxUpdate_3[3:0]) begin
            TBEValid_14 <= 1'h0;
          end else begin
            TBEValid_14 <= _GEN_1539;
          end
        end else begin
          TBEValid_14 <= _GEN_1539;
        end
      end else if (isAlloc_5) begin
        TBEValid_14 <= _GEN_2648;
      end else if (_T_199) begin
        if (4'he == idxUpdate_5[3:0]) begin
          TBEValid_14 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_14 <= _GEN_2134;
        end else if (_T_177) begin
          if (4'he == idxUpdate_4[3:0]) begin
            TBEValid_14 <= 1'h0;
          end else begin
            TBEValid_14 <= _GEN_2053;
          end
        end else begin
          TBEValid_14 <= _GEN_2053;
        end
      end else if (isAlloc_4) begin
        TBEValid_14 <= _GEN_2134;
      end else if (_T_177) begin
        if (4'he == idxUpdate_4[3:0]) begin
          TBEValid_14 <= 1'h0;
        end else begin
          TBEValid_14 <= _GEN_2053;
        end
      end else begin
        TBEValid_14 <= _GEN_2053;
      end
    end else if (isAlloc_6) begin
      TBEValid_14 <= _GEN_3162;
    end else if (_T_221) begin
      if (4'he == idxUpdate_6[3:0]) begin
        TBEValid_14 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_14 <= _GEN_2648;
      end else if (_T_199) begin
        if (4'he == idxUpdate_5[3:0]) begin
          TBEValid_14 <= 1'h0;
        end else begin
          TBEValid_14 <= _GEN_2567;
        end
      end else begin
        TBEValid_14 <= _GEN_2567;
      end
    end else if (isAlloc_5) begin
      TBEValid_14 <= _GEN_2648;
    end else if (_T_199) begin
      if (4'he == idxUpdate_5[3:0]) begin
        TBEValid_14 <= 1'h0;
      end else begin
        TBEValid_14 <= _GEN_2567;
      end
    end else begin
      TBEValid_14 <= _GEN_2567;
    end
    if (reset) begin
      TBEValid_15 <= 1'h0;
    end else if (isAlloc_7) begin
      TBEValid_15 <= _GEN_3677;
    end else if (_T_243) begin
      if (4'hf == idxUpdate_7[3:0]) begin
        TBEValid_15 <= 1'h0;
      end else if (isAlloc_6) begin
        TBEValid_15 <= _GEN_3163;
      end else if (_T_221) begin
        if (4'hf == idxUpdate_6[3:0]) begin
          TBEValid_15 <= 1'h0;
        end else if (isAlloc_5) begin
          TBEValid_15 <= _GEN_2649;
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEValid_15 <= 1'h0;
          end else if (isAlloc_4) begin
            TBEValid_15 <= _GEN_2135;
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEValid_15 <= 1'h0;
            end else if (isAlloc_3) begin
              TBEValid_15 <= _GEN_1621;
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEValid_15 <= 1'h0;
              end else if (isAlloc_2) begin
                TBEValid_15 <= _GEN_1107;
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEValid_15 <= 1'h0;
                end else if (isAlloc_1) begin
                  TBEValid_15 <= _GEN_593;
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEValid_15 <= 1'h0;
                  end else if (isAlloc_0) begin
                    TBEValid_15 <= _GEN_79;
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEValid_15 <= 1'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  TBEValid_15 <= _GEN_79;
                end else if (_T_89) begin
                  if (4'hf == idxUpdate_0[3:0]) begin
                    TBEValid_15 <= 1'h0;
                  end
                end
              end else if (isAlloc_1) begin
                TBEValid_15 <= _GEN_593;
              end else if (_T_111) begin
                if (4'hf == idxUpdate_1[3:0]) begin
                  TBEValid_15 <= 1'h0;
                end else if (isAlloc_0) begin
                  TBEValid_15 <= _GEN_79;
                end else if (_T_89) begin
                  if (4'hf == idxUpdate_0[3:0]) begin
                    TBEValid_15 <= 1'h0;
                  end
                end
              end else if (isAlloc_0) begin
                TBEValid_15 <= _GEN_79;
              end else if (_T_89) begin
                if (4'hf == idxUpdate_0[3:0]) begin
                  TBEValid_15 <= 1'h0;
                end
              end
            end else if (isAlloc_2) begin
              TBEValid_15 <= _GEN_1107;
            end else if (_T_133) begin
              if (4'hf == idxUpdate_2[3:0]) begin
                TBEValid_15 <= 1'h0;
              end else if (isAlloc_1) begin
                TBEValid_15 <= _GEN_593;
              end else if (_T_111) begin
                if (4'hf == idxUpdate_1[3:0]) begin
                  TBEValid_15 <= 1'h0;
                end else begin
                  TBEValid_15 <= _GEN_512;
                end
              end else begin
                TBEValid_15 <= _GEN_512;
              end
            end else if (isAlloc_1) begin
              TBEValid_15 <= _GEN_593;
            end else if (_T_111) begin
              if (4'hf == idxUpdate_1[3:0]) begin
                TBEValid_15 <= 1'h0;
              end else begin
                TBEValid_15 <= _GEN_512;
              end
            end else begin
              TBEValid_15 <= _GEN_512;
            end
          end else if (isAlloc_3) begin
            TBEValid_15 <= _GEN_1621;
          end else if (_T_155) begin
            if (4'hf == idxUpdate_3[3:0]) begin
              TBEValid_15 <= 1'h0;
            end else if (isAlloc_2) begin
              TBEValid_15 <= _GEN_1107;
            end else if (_T_133) begin
              if (4'hf == idxUpdate_2[3:0]) begin
                TBEValid_15 <= 1'h0;
              end else begin
                TBEValid_15 <= _GEN_1026;
              end
            end else begin
              TBEValid_15 <= _GEN_1026;
            end
          end else if (isAlloc_2) begin
            TBEValid_15 <= _GEN_1107;
          end else if (_T_133) begin
            if (4'hf == idxUpdate_2[3:0]) begin
              TBEValid_15 <= 1'h0;
            end else begin
              TBEValid_15 <= _GEN_1026;
            end
          end else begin
            TBEValid_15 <= _GEN_1026;
          end
        end else if (isAlloc_4) begin
          TBEValid_15 <= _GEN_2135;
        end else if (_T_177) begin
          if (4'hf == idxUpdate_4[3:0]) begin
            TBEValid_15 <= 1'h0;
          end else if (isAlloc_3) begin
            TBEValid_15 <= _GEN_1621;
          end else if (_T_155) begin
            if (4'hf == idxUpdate_3[3:0]) begin
              TBEValid_15 <= 1'h0;
            end else begin
              TBEValid_15 <= _GEN_1540;
            end
          end else begin
            TBEValid_15 <= _GEN_1540;
          end
        end else if (isAlloc_3) begin
          TBEValid_15 <= _GEN_1621;
        end else if (_T_155) begin
          if (4'hf == idxUpdate_3[3:0]) begin
            TBEValid_15 <= 1'h0;
          end else begin
            TBEValid_15 <= _GEN_1540;
          end
        end else begin
          TBEValid_15 <= _GEN_1540;
        end
      end else if (isAlloc_5) begin
        TBEValid_15 <= _GEN_2649;
      end else if (_T_199) begin
        if (4'hf == idxUpdate_5[3:0]) begin
          TBEValid_15 <= 1'h0;
        end else if (isAlloc_4) begin
          TBEValid_15 <= _GEN_2135;
        end else if (_T_177) begin
          if (4'hf == idxUpdate_4[3:0]) begin
            TBEValid_15 <= 1'h0;
          end else begin
            TBEValid_15 <= _GEN_2054;
          end
        end else begin
          TBEValid_15 <= _GEN_2054;
        end
      end else if (isAlloc_4) begin
        TBEValid_15 <= _GEN_2135;
      end else if (_T_177) begin
        if (4'hf == idxUpdate_4[3:0]) begin
          TBEValid_15 <= 1'h0;
        end else begin
          TBEValid_15 <= _GEN_2054;
        end
      end else begin
        TBEValid_15 <= _GEN_2054;
      end
    end else if (isAlloc_6) begin
      TBEValid_15 <= _GEN_3163;
    end else if (_T_221) begin
      if (4'hf == idxUpdate_6[3:0]) begin
        TBEValid_15 <= 1'h0;
      end else if (isAlloc_5) begin
        TBEValid_15 <= _GEN_2649;
      end else if (_T_199) begin
        if (4'hf == idxUpdate_5[3:0]) begin
          TBEValid_15 <= 1'h0;
        end else begin
          TBEValid_15 <= _GEN_2568;
        end
      end else begin
        TBEValid_15 <= _GEN_2568;
      end
    end else if (isAlloc_5) begin
      TBEValid_15 <= _GEN_2649;
    end else if (_T_199) begin
      if (4'hf == idxUpdate_5[3:0]) begin
        TBEValid_15 <= 1'h0;
      end else begin
        TBEValid_15 <= _GEN_2568;
      end
    end else begin
      TBEValid_15 <= _GEN_2568;
    end
    if (reset) begin
      TBEAddr_0 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h0 == idxAlloc[3:0]) begin
        TBEAddr_0 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'h0 == idxAlloc[3:0]) begin
          TBEAddr_0 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEAddr_0 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEAddr_0 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEAddr_0 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEAddr_0 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEAddr_0 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEAddr_0 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEAddr_0 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEAddr_0 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEAddr_0 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEAddr_0 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEAddr_0 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'h0 == idxUpdate_0[3:0]) begin
                    TBEAddr_0 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEAddr_0 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEAddr_0 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h0 == idxAlloc[3:0]) begin
                      TBEAddr_0 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h0 == idxUpdate_0[3:0]) begin
                      TBEAddr_0 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEAddr_0 <= 32'h0;
                  end else begin
                    TBEAddr_0 <= _GEN_481;
                  end
                end else begin
                  TBEAddr_0 <= _GEN_481;
                end
              end else if (isAlloc_1) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEAddr_0 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_0 <= _GEN_481;
                end
              end else if (_T_111) begin
                if (4'h0 == idxUpdate_1[3:0]) begin
                  TBEAddr_0 <= 32'h0;
                end else begin
                  TBEAddr_0 <= _GEN_481;
                end
              end else begin
                TBEAddr_0 <= _GEN_481;
              end
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEAddr_0 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEAddr_0 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h0 == idxAlloc[3:0]) begin
                    TBEAddr_0 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_0 <= _GEN_481;
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUpdate_1[3:0]) begin
                    TBEAddr_0 <= 32'h0;
                  end else begin
                    TBEAddr_0 <= _GEN_481;
                  end
                end else begin
                  TBEAddr_0 <= _GEN_481;
                end
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEAddr_0 <= 32'h0;
                end else begin
                  TBEAddr_0 <= _GEN_995;
                end
              end else begin
                TBEAddr_0 <= _GEN_995;
              end
            end else if (isAlloc_2) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEAddr_0 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_0 <= _GEN_995;
              end
            end else if (_T_133) begin
              if (4'h0 == idxUpdate_2[3:0]) begin
                TBEAddr_0 <= 32'h0;
              end else begin
                TBEAddr_0 <= _GEN_995;
              end
            end else begin
              TBEAddr_0 <= _GEN_995;
            end
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEAddr_0 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEAddr_0 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h0 == idxAlloc[3:0]) begin
                  TBEAddr_0 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_0 <= _GEN_995;
                end
              end else if (_T_133) begin
                if (4'h0 == idxUpdate_2[3:0]) begin
                  TBEAddr_0 <= 32'h0;
                end else begin
                  TBEAddr_0 <= _GEN_995;
                end
              end else begin
                TBEAddr_0 <= _GEN_995;
              end
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEAddr_0 <= 32'h0;
              end else begin
                TBEAddr_0 <= _GEN_1509;
              end
            end else begin
              TBEAddr_0 <= _GEN_1509;
            end
          end else if (isAlloc_3) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEAddr_0 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_0 <= _GEN_1509;
            end
          end else if (_T_155) begin
            if (4'h0 == idxUpdate_3[3:0]) begin
              TBEAddr_0 <= 32'h0;
            end else begin
              TBEAddr_0 <= _GEN_1509;
            end
          end else begin
            TBEAddr_0 <= _GEN_1509;
          end
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEAddr_0 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEAddr_0 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h0 == idxAlloc[3:0]) begin
                TBEAddr_0 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_0 <= _GEN_1509;
              end
            end else if (_T_155) begin
              if (4'h0 == idxUpdate_3[3:0]) begin
                TBEAddr_0 <= 32'h0;
              end else begin
                TBEAddr_0 <= _GEN_1509;
              end
            end else begin
              TBEAddr_0 <= _GEN_1509;
            end
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEAddr_0 <= 32'h0;
            end else begin
              TBEAddr_0 <= _GEN_2023;
            end
          end else begin
            TBEAddr_0 <= _GEN_2023;
          end
        end else if (isAlloc_4) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEAddr_0 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_0 <= _GEN_2023;
          end
        end else if (_T_177) begin
          if (4'h0 == idxUpdate_4[3:0]) begin
            TBEAddr_0 <= 32'h0;
          end else begin
            TBEAddr_0 <= _GEN_2023;
          end
        end else begin
          TBEAddr_0 <= _GEN_2023;
        end
      end else if (_T_221) begin
        if (4'h0 == idxUpdate_6[3:0]) begin
          TBEAddr_0 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEAddr_0 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h0 == idxAlloc[3:0]) begin
              TBEAddr_0 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_0 <= _GEN_2023;
            end
          end else if (_T_177) begin
            if (4'h0 == idxUpdate_4[3:0]) begin
              TBEAddr_0 <= 32'h0;
            end else begin
              TBEAddr_0 <= _GEN_2023;
            end
          end else begin
            TBEAddr_0 <= _GEN_2023;
          end
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEAddr_0 <= 32'h0;
          end else begin
            TBEAddr_0 <= _GEN_2537;
          end
        end else begin
          TBEAddr_0 <= _GEN_2537;
        end
      end else if (isAlloc_5) begin
        if (4'h0 == idxAlloc[3:0]) begin
          TBEAddr_0 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_0 <= _GEN_2537;
        end
      end else if (_T_199) begin
        if (4'h0 == idxUpdate_5[3:0]) begin
          TBEAddr_0 <= 32'h0;
        end else begin
          TBEAddr_0 <= _GEN_2537;
        end
      end else begin
        TBEAddr_0 <= _GEN_2537;
      end
    end else if (_T_243) begin
      if (4'h0 == idxUpdate_7[3:0]) begin
        TBEAddr_0 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h0 == idxAlloc[3:0]) begin
          TBEAddr_0 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h0 == idxAlloc[3:0]) begin
            TBEAddr_0 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_0 <= _GEN_2537;
          end
        end else if (_T_199) begin
          if (4'h0 == idxUpdate_5[3:0]) begin
            TBEAddr_0 <= 32'h0;
          end else begin
            TBEAddr_0 <= _GEN_2537;
          end
        end else begin
          TBEAddr_0 <= _GEN_2537;
        end
      end else if (_T_221) begin
        if (4'h0 == idxUpdate_6[3:0]) begin
          TBEAddr_0 <= 32'h0;
        end else begin
          TBEAddr_0 <= _GEN_3051;
        end
      end else begin
        TBEAddr_0 <= _GEN_3051;
      end
    end else if (isAlloc_6) begin
      if (4'h0 == idxAlloc[3:0]) begin
        TBEAddr_0 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_0 <= _GEN_3051;
      end
    end else if (_T_221) begin
      if (4'h0 == idxUpdate_6[3:0]) begin
        TBEAddr_0 <= 32'h0;
      end else begin
        TBEAddr_0 <= _GEN_3051;
      end
    end else begin
      TBEAddr_0 <= _GEN_3051;
    end
    if (reset) begin
      TBEAddr_1 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h1 == idxAlloc[3:0]) begin
        TBEAddr_1 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'h1 == idxAlloc[3:0]) begin
          TBEAddr_1 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEAddr_1 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEAddr_1 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEAddr_1 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEAddr_1 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEAddr_1 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEAddr_1 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEAddr_1 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEAddr_1 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEAddr_1 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEAddr_1 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEAddr_1 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'h1 == idxUpdate_0[3:0]) begin
                    TBEAddr_1 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEAddr_1 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEAddr_1 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h1 == idxAlloc[3:0]) begin
                      TBEAddr_1 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h1 == idxUpdate_0[3:0]) begin
                      TBEAddr_1 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEAddr_1 <= 32'h0;
                  end else begin
                    TBEAddr_1 <= _GEN_482;
                  end
                end else begin
                  TBEAddr_1 <= _GEN_482;
                end
              end else if (isAlloc_1) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEAddr_1 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_1 <= _GEN_482;
                end
              end else if (_T_111) begin
                if (4'h1 == idxUpdate_1[3:0]) begin
                  TBEAddr_1 <= 32'h0;
                end else begin
                  TBEAddr_1 <= _GEN_482;
                end
              end else begin
                TBEAddr_1 <= _GEN_482;
              end
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEAddr_1 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEAddr_1 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h1 == idxAlloc[3:0]) begin
                    TBEAddr_1 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_1 <= _GEN_482;
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUpdate_1[3:0]) begin
                    TBEAddr_1 <= 32'h0;
                  end else begin
                    TBEAddr_1 <= _GEN_482;
                  end
                end else begin
                  TBEAddr_1 <= _GEN_482;
                end
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEAddr_1 <= 32'h0;
                end else begin
                  TBEAddr_1 <= _GEN_996;
                end
              end else begin
                TBEAddr_1 <= _GEN_996;
              end
            end else if (isAlloc_2) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEAddr_1 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_1 <= _GEN_996;
              end
            end else if (_T_133) begin
              if (4'h1 == idxUpdate_2[3:0]) begin
                TBEAddr_1 <= 32'h0;
              end else begin
                TBEAddr_1 <= _GEN_996;
              end
            end else begin
              TBEAddr_1 <= _GEN_996;
            end
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEAddr_1 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEAddr_1 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h1 == idxAlloc[3:0]) begin
                  TBEAddr_1 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_1 <= _GEN_996;
                end
              end else if (_T_133) begin
                if (4'h1 == idxUpdate_2[3:0]) begin
                  TBEAddr_1 <= 32'h0;
                end else begin
                  TBEAddr_1 <= _GEN_996;
                end
              end else begin
                TBEAddr_1 <= _GEN_996;
              end
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEAddr_1 <= 32'h0;
              end else begin
                TBEAddr_1 <= _GEN_1510;
              end
            end else begin
              TBEAddr_1 <= _GEN_1510;
            end
          end else if (isAlloc_3) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEAddr_1 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_1 <= _GEN_1510;
            end
          end else if (_T_155) begin
            if (4'h1 == idxUpdate_3[3:0]) begin
              TBEAddr_1 <= 32'h0;
            end else begin
              TBEAddr_1 <= _GEN_1510;
            end
          end else begin
            TBEAddr_1 <= _GEN_1510;
          end
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEAddr_1 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEAddr_1 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h1 == idxAlloc[3:0]) begin
                TBEAddr_1 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_1 <= _GEN_1510;
              end
            end else if (_T_155) begin
              if (4'h1 == idxUpdate_3[3:0]) begin
                TBEAddr_1 <= 32'h0;
              end else begin
                TBEAddr_1 <= _GEN_1510;
              end
            end else begin
              TBEAddr_1 <= _GEN_1510;
            end
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEAddr_1 <= 32'h0;
            end else begin
              TBEAddr_1 <= _GEN_2024;
            end
          end else begin
            TBEAddr_1 <= _GEN_2024;
          end
        end else if (isAlloc_4) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEAddr_1 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_1 <= _GEN_2024;
          end
        end else if (_T_177) begin
          if (4'h1 == idxUpdate_4[3:0]) begin
            TBEAddr_1 <= 32'h0;
          end else begin
            TBEAddr_1 <= _GEN_2024;
          end
        end else begin
          TBEAddr_1 <= _GEN_2024;
        end
      end else if (_T_221) begin
        if (4'h1 == idxUpdate_6[3:0]) begin
          TBEAddr_1 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEAddr_1 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h1 == idxAlloc[3:0]) begin
              TBEAddr_1 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_1 <= _GEN_2024;
            end
          end else if (_T_177) begin
            if (4'h1 == idxUpdate_4[3:0]) begin
              TBEAddr_1 <= 32'h0;
            end else begin
              TBEAddr_1 <= _GEN_2024;
            end
          end else begin
            TBEAddr_1 <= _GEN_2024;
          end
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEAddr_1 <= 32'h0;
          end else begin
            TBEAddr_1 <= _GEN_2538;
          end
        end else begin
          TBEAddr_1 <= _GEN_2538;
        end
      end else if (isAlloc_5) begin
        if (4'h1 == idxAlloc[3:0]) begin
          TBEAddr_1 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_1 <= _GEN_2538;
        end
      end else if (_T_199) begin
        if (4'h1 == idxUpdate_5[3:0]) begin
          TBEAddr_1 <= 32'h0;
        end else begin
          TBEAddr_1 <= _GEN_2538;
        end
      end else begin
        TBEAddr_1 <= _GEN_2538;
      end
    end else if (_T_243) begin
      if (4'h1 == idxUpdate_7[3:0]) begin
        TBEAddr_1 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h1 == idxAlloc[3:0]) begin
          TBEAddr_1 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h1 == idxAlloc[3:0]) begin
            TBEAddr_1 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_1 <= _GEN_2538;
          end
        end else if (_T_199) begin
          if (4'h1 == idxUpdate_5[3:0]) begin
            TBEAddr_1 <= 32'h0;
          end else begin
            TBEAddr_1 <= _GEN_2538;
          end
        end else begin
          TBEAddr_1 <= _GEN_2538;
        end
      end else if (_T_221) begin
        if (4'h1 == idxUpdate_6[3:0]) begin
          TBEAddr_1 <= 32'h0;
        end else begin
          TBEAddr_1 <= _GEN_3052;
        end
      end else begin
        TBEAddr_1 <= _GEN_3052;
      end
    end else if (isAlloc_6) begin
      if (4'h1 == idxAlloc[3:0]) begin
        TBEAddr_1 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_1 <= _GEN_3052;
      end
    end else if (_T_221) begin
      if (4'h1 == idxUpdate_6[3:0]) begin
        TBEAddr_1 <= 32'h0;
      end else begin
        TBEAddr_1 <= _GEN_3052;
      end
    end else begin
      TBEAddr_1 <= _GEN_3052;
    end
    if (reset) begin
      TBEAddr_2 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h2 == idxAlloc[3:0]) begin
        TBEAddr_2 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'h2 == idxAlloc[3:0]) begin
          TBEAddr_2 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEAddr_2 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEAddr_2 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEAddr_2 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEAddr_2 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEAddr_2 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEAddr_2 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEAddr_2 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEAddr_2 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEAddr_2 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEAddr_2 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEAddr_2 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'h2 == idxUpdate_0[3:0]) begin
                    TBEAddr_2 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEAddr_2 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEAddr_2 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h2 == idxAlloc[3:0]) begin
                      TBEAddr_2 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h2 == idxUpdate_0[3:0]) begin
                      TBEAddr_2 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEAddr_2 <= 32'h0;
                  end else begin
                    TBEAddr_2 <= _GEN_483;
                  end
                end else begin
                  TBEAddr_2 <= _GEN_483;
                end
              end else if (isAlloc_1) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEAddr_2 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_2 <= _GEN_483;
                end
              end else if (_T_111) begin
                if (4'h2 == idxUpdate_1[3:0]) begin
                  TBEAddr_2 <= 32'h0;
                end else begin
                  TBEAddr_2 <= _GEN_483;
                end
              end else begin
                TBEAddr_2 <= _GEN_483;
              end
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEAddr_2 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEAddr_2 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h2 == idxAlloc[3:0]) begin
                    TBEAddr_2 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_2 <= _GEN_483;
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUpdate_1[3:0]) begin
                    TBEAddr_2 <= 32'h0;
                  end else begin
                    TBEAddr_2 <= _GEN_483;
                  end
                end else begin
                  TBEAddr_2 <= _GEN_483;
                end
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEAddr_2 <= 32'h0;
                end else begin
                  TBEAddr_2 <= _GEN_997;
                end
              end else begin
                TBEAddr_2 <= _GEN_997;
              end
            end else if (isAlloc_2) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEAddr_2 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_2 <= _GEN_997;
              end
            end else if (_T_133) begin
              if (4'h2 == idxUpdate_2[3:0]) begin
                TBEAddr_2 <= 32'h0;
              end else begin
                TBEAddr_2 <= _GEN_997;
              end
            end else begin
              TBEAddr_2 <= _GEN_997;
            end
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEAddr_2 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEAddr_2 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h2 == idxAlloc[3:0]) begin
                  TBEAddr_2 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_2 <= _GEN_997;
                end
              end else if (_T_133) begin
                if (4'h2 == idxUpdate_2[3:0]) begin
                  TBEAddr_2 <= 32'h0;
                end else begin
                  TBEAddr_2 <= _GEN_997;
                end
              end else begin
                TBEAddr_2 <= _GEN_997;
              end
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEAddr_2 <= 32'h0;
              end else begin
                TBEAddr_2 <= _GEN_1511;
              end
            end else begin
              TBEAddr_2 <= _GEN_1511;
            end
          end else if (isAlloc_3) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEAddr_2 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_2 <= _GEN_1511;
            end
          end else if (_T_155) begin
            if (4'h2 == idxUpdate_3[3:0]) begin
              TBEAddr_2 <= 32'h0;
            end else begin
              TBEAddr_2 <= _GEN_1511;
            end
          end else begin
            TBEAddr_2 <= _GEN_1511;
          end
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEAddr_2 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEAddr_2 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h2 == idxAlloc[3:0]) begin
                TBEAddr_2 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_2 <= _GEN_1511;
              end
            end else if (_T_155) begin
              if (4'h2 == idxUpdate_3[3:0]) begin
                TBEAddr_2 <= 32'h0;
              end else begin
                TBEAddr_2 <= _GEN_1511;
              end
            end else begin
              TBEAddr_2 <= _GEN_1511;
            end
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEAddr_2 <= 32'h0;
            end else begin
              TBEAddr_2 <= _GEN_2025;
            end
          end else begin
            TBEAddr_2 <= _GEN_2025;
          end
        end else if (isAlloc_4) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEAddr_2 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_2 <= _GEN_2025;
          end
        end else if (_T_177) begin
          if (4'h2 == idxUpdate_4[3:0]) begin
            TBEAddr_2 <= 32'h0;
          end else begin
            TBEAddr_2 <= _GEN_2025;
          end
        end else begin
          TBEAddr_2 <= _GEN_2025;
        end
      end else if (_T_221) begin
        if (4'h2 == idxUpdate_6[3:0]) begin
          TBEAddr_2 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEAddr_2 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h2 == idxAlloc[3:0]) begin
              TBEAddr_2 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_2 <= _GEN_2025;
            end
          end else if (_T_177) begin
            if (4'h2 == idxUpdate_4[3:0]) begin
              TBEAddr_2 <= 32'h0;
            end else begin
              TBEAddr_2 <= _GEN_2025;
            end
          end else begin
            TBEAddr_2 <= _GEN_2025;
          end
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEAddr_2 <= 32'h0;
          end else begin
            TBEAddr_2 <= _GEN_2539;
          end
        end else begin
          TBEAddr_2 <= _GEN_2539;
        end
      end else if (isAlloc_5) begin
        if (4'h2 == idxAlloc[3:0]) begin
          TBEAddr_2 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_2 <= _GEN_2539;
        end
      end else if (_T_199) begin
        if (4'h2 == idxUpdate_5[3:0]) begin
          TBEAddr_2 <= 32'h0;
        end else begin
          TBEAddr_2 <= _GEN_2539;
        end
      end else begin
        TBEAddr_2 <= _GEN_2539;
      end
    end else if (_T_243) begin
      if (4'h2 == idxUpdate_7[3:0]) begin
        TBEAddr_2 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h2 == idxAlloc[3:0]) begin
          TBEAddr_2 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h2 == idxAlloc[3:0]) begin
            TBEAddr_2 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_2 <= _GEN_2539;
          end
        end else if (_T_199) begin
          if (4'h2 == idxUpdate_5[3:0]) begin
            TBEAddr_2 <= 32'h0;
          end else begin
            TBEAddr_2 <= _GEN_2539;
          end
        end else begin
          TBEAddr_2 <= _GEN_2539;
        end
      end else if (_T_221) begin
        if (4'h2 == idxUpdate_6[3:0]) begin
          TBEAddr_2 <= 32'h0;
        end else begin
          TBEAddr_2 <= _GEN_3053;
        end
      end else begin
        TBEAddr_2 <= _GEN_3053;
      end
    end else if (isAlloc_6) begin
      if (4'h2 == idxAlloc[3:0]) begin
        TBEAddr_2 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_2 <= _GEN_3053;
      end
    end else if (_T_221) begin
      if (4'h2 == idxUpdate_6[3:0]) begin
        TBEAddr_2 <= 32'h0;
      end else begin
        TBEAddr_2 <= _GEN_3053;
      end
    end else begin
      TBEAddr_2 <= _GEN_3053;
    end
    if (reset) begin
      TBEAddr_3 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h3 == idxAlloc[3:0]) begin
        TBEAddr_3 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'h3 == idxAlloc[3:0]) begin
          TBEAddr_3 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEAddr_3 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEAddr_3 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEAddr_3 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEAddr_3 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEAddr_3 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEAddr_3 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEAddr_3 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEAddr_3 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEAddr_3 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEAddr_3 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEAddr_3 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'h3 == idxUpdate_0[3:0]) begin
                    TBEAddr_3 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEAddr_3 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEAddr_3 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h3 == idxAlloc[3:0]) begin
                      TBEAddr_3 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h3 == idxUpdate_0[3:0]) begin
                      TBEAddr_3 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEAddr_3 <= 32'h0;
                  end else begin
                    TBEAddr_3 <= _GEN_484;
                  end
                end else begin
                  TBEAddr_3 <= _GEN_484;
                end
              end else if (isAlloc_1) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEAddr_3 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_3 <= _GEN_484;
                end
              end else if (_T_111) begin
                if (4'h3 == idxUpdate_1[3:0]) begin
                  TBEAddr_3 <= 32'h0;
                end else begin
                  TBEAddr_3 <= _GEN_484;
                end
              end else begin
                TBEAddr_3 <= _GEN_484;
              end
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEAddr_3 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEAddr_3 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h3 == idxAlloc[3:0]) begin
                    TBEAddr_3 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_3 <= _GEN_484;
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUpdate_1[3:0]) begin
                    TBEAddr_3 <= 32'h0;
                  end else begin
                    TBEAddr_3 <= _GEN_484;
                  end
                end else begin
                  TBEAddr_3 <= _GEN_484;
                end
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEAddr_3 <= 32'h0;
                end else begin
                  TBEAddr_3 <= _GEN_998;
                end
              end else begin
                TBEAddr_3 <= _GEN_998;
              end
            end else if (isAlloc_2) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEAddr_3 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_3 <= _GEN_998;
              end
            end else if (_T_133) begin
              if (4'h3 == idxUpdate_2[3:0]) begin
                TBEAddr_3 <= 32'h0;
              end else begin
                TBEAddr_3 <= _GEN_998;
              end
            end else begin
              TBEAddr_3 <= _GEN_998;
            end
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEAddr_3 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEAddr_3 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h3 == idxAlloc[3:0]) begin
                  TBEAddr_3 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_3 <= _GEN_998;
                end
              end else if (_T_133) begin
                if (4'h3 == idxUpdate_2[3:0]) begin
                  TBEAddr_3 <= 32'h0;
                end else begin
                  TBEAddr_3 <= _GEN_998;
                end
              end else begin
                TBEAddr_3 <= _GEN_998;
              end
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEAddr_3 <= 32'h0;
              end else begin
                TBEAddr_3 <= _GEN_1512;
              end
            end else begin
              TBEAddr_3 <= _GEN_1512;
            end
          end else if (isAlloc_3) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEAddr_3 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_3 <= _GEN_1512;
            end
          end else if (_T_155) begin
            if (4'h3 == idxUpdate_3[3:0]) begin
              TBEAddr_3 <= 32'h0;
            end else begin
              TBEAddr_3 <= _GEN_1512;
            end
          end else begin
            TBEAddr_3 <= _GEN_1512;
          end
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEAddr_3 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEAddr_3 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h3 == idxAlloc[3:0]) begin
                TBEAddr_3 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_3 <= _GEN_1512;
              end
            end else if (_T_155) begin
              if (4'h3 == idxUpdate_3[3:0]) begin
                TBEAddr_3 <= 32'h0;
              end else begin
                TBEAddr_3 <= _GEN_1512;
              end
            end else begin
              TBEAddr_3 <= _GEN_1512;
            end
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEAddr_3 <= 32'h0;
            end else begin
              TBEAddr_3 <= _GEN_2026;
            end
          end else begin
            TBEAddr_3 <= _GEN_2026;
          end
        end else if (isAlloc_4) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEAddr_3 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_3 <= _GEN_2026;
          end
        end else if (_T_177) begin
          if (4'h3 == idxUpdate_4[3:0]) begin
            TBEAddr_3 <= 32'h0;
          end else begin
            TBEAddr_3 <= _GEN_2026;
          end
        end else begin
          TBEAddr_3 <= _GEN_2026;
        end
      end else if (_T_221) begin
        if (4'h3 == idxUpdate_6[3:0]) begin
          TBEAddr_3 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEAddr_3 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h3 == idxAlloc[3:0]) begin
              TBEAddr_3 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_3 <= _GEN_2026;
            end
          end else if (_T_177) begin
            if (4'h3 == idxUpdate_4[3:0]) begin
              TBEAddr_3 <= 32'h0;
            end else begin
              TBEAddr_3 <= _GEN_2026;
            end
          end else begin
            TBEAddr_3 <= _GEN_2026;
          end
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEAddr_3 <= 32'h0;
          end else begin
            TBEAddr_3 <= _GEN_2540;
          end
        end else begin
          TBEAddr_3 <= _GEN_2540;
        end
      end else if (isAlloc_5) begin
        if (4'h3 == idxAlloc[3:0]) begin
          TBEAddr_3 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_3 <= _GEN_2540;
        end
      end else if (_T_199) begin
        if (4'h3 == idxUpdate_5[3:0]) begin
          TBEAddr_3 <= 32'h0;
        end else begin
          TBEAddr_3 <= _GEN_2540;
        end
      end else begin
        TBEAddr_3 <= _GEN_2540;
      end
    end else if (_T_243) begin
      if (4'h3 == idxUpdate_7[3:0]) begin
        TBEAddr_3 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h3 == idxAlloc[3:0]) begin
          TBEAddr_3 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h3 == idxAlloc[3:0]) begin
            TBEAddr_3 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_3 <= _GEN_2540;
          end
        end else if (_T_199) begin
          if (4'h3 == idxUpdate_5[3:0]) begin
            TBEAddr_3 <= 32'h0;
          end else begin
            TBEAddr_3 <= _GEN_2540;
          end
        end else begin
          TBEAddr_3 <= _GEN_2540;
        end
      end else if (_T_221) begin
        if (4'h3 == idxUpdate_6[3:0]) begin
          TBEAddr_3 <= 32'h0;
        end else begin
          TBEAddr_3 <= _GEN_3054;
        end
      end else begin
        TBEAddr_3 <= _GEN_3054;
      end
    end else if (isAlloc_6) begin
      if (4'h3 == idxAlloc[3:0]) begin
        TBEAddr_3 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_3 <= _GEN_3054;
      end
    end else if (_T_221) begin
      if (4'h3 == idxUpdate_6[3:0]) begin
        TBEAddr_3 <= 32'h0;
      end else begin
        TBEAddr_3 <= _GEN_3054;
      end
    end else begin
      TBEAddr_3 <= _GEN_3054;
    end
    if (reset) begin
      TBEAddr_4 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h4 == idxAlloc[3:0]) begin
        TBEAddr_4 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'h4 == idxAlloc[3:0]) begin
          TBEAddr_4 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEAddr_4 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEAddr_4 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEAddr_4 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEAddr_4 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEAddr_4 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEAddr_4 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEAddr_4 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEAddr_4 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEAddr_4 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEAddr_4 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEAddr_4 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'h4 == idxUpdate_0[3:0]) begin
                    TBEAddr_4 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEAddr_4 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEAddr_4 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h4 == idxAlloc[3:0]) begin
                      TBEAddr_4 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h4 == idxUpdate_0[3:0]) begin
                      TBEAddr_4 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEAddr_4 <= 32'h0;
                  end else begin
                    TBEAddr_4 <= _GEN_485;
                  end
                end else begin
                  TBEAddr_4 <= _GEN_485;
                end
              end else if (isAlloc_1) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEAddr_4 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_4 <= _GEN_485;
                end
              end else if (_T_111) begin
                if (4'h4 == idxUpdate_1[3:0]) begin
                  TBEAddr_4 <= 32'h0;
                end else begin
                  TBEAddr_4 <= _GEN_485;
                end
              end else begin
                TBEAddr_4 <= _GEN_485;
              end
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEAddr_4 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEAddr_4 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h4 == idxAlloc[3:0]) begin
                    TBEAddr_4 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_4 <= _GEN_485;
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUpdate_1[3:0]) begin
                    TBEAddr_4 <= 32'h0;
                  end else begin
                    TBEAddr_4 <= _GEN_485;
                  end
                end else begin
                  TBEAddr_4 <= _GEN_485;
                end
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEAddr_4 <= 32'h0;
                end else begin
                  TBEAddr_4 <= _GEN_999;
                end
              end else begin
                TBEAddr_4 <= _GEN_999;
              end
            end else if (isAlloc_2) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEAddr_4 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_4 <= _GEN_999;
              end
            end else if (_T_133) begin
              if (4'h4 == idxUpdate_2[3:0]) begin
                TBEAddr_4 <= 32'h0;
              end else begin
                TBEAddr_4 <= _GEN_999;
              end
            end else begin
              TBEAddr_4 <= _GEN_999;
            end
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEAddr_4 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEAddr_4 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h4 == idxAlloc[3:0]) begin
                  TBEAddr_4 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_4 <= _GEN_999;
                end
              end else if (_T_133) begin
                if (4'h4 == idxUpdate_2[3:0]) begin
                  TBEAddr_4 <= 32'h0;
                end else begin
                  TBEAddr_4 <= _GEN_999;
                end
              end else begin
                TBEAddr_4 <= _GEN_999;
              end
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEAddr_4 <= 32'h0;
              end else begin
                TBEAddr_4 <= _GEN_1513;
              end
            end else begin
              TBEAddr_4 <= _GEN_1513;
            end
          end else if (isAlloc_3) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEAddr_4 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_4 <= _GEN_1513;
            end
          end else if (_T_155) begin
            if (4'h4 == idxUpdate_3[3:0]) begin
              TBEAddr_4 <= 32'h0;
            end else begin
              TBEAddr_4 <= _GEN_1513;
            end
          end else begin
            TBEAddr_4 <= _GEN_1513;
          end
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEAddr_4 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEAddr_4 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h4 == idxAlloc[3:0]) begin
                TBEAddr_4 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_4 <= _GEN_1513;
              end
            end else if (_T_155) begin
              if (4'h4 == idxUpdate_3[3:0]) begin
                TBEAddr_4 <= 32'h0;
              end else begin
                TBEAddr_4 <= _GEN_1513;
              end
            end else begin
              TBEAddr_4 <= _GEN_1513;
            end
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEAddr_4 <= 32'h0;
            end else begin
              TBEAddr_4 <= _GEN_2027;
            end
          end else begin
            TBEAddr_4 <= _GEN_2027;
          end
        end else if (isAlloc_4) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEAddr_4 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_4 <= _GEN_2027;
          end
        end else if (_T_177) begin
          if (4'h4 == idxUpdate_4[3:0]) begin
            TBEAddr_4 <= 32'h0;
          end else begin
            TBEAddr_4 <= _GEN_2027;
          end
        end else begin
          TBEAddr_4 <= _GEN_2027;
        end
      end else if (_T_221) begin
        if (4'h4 == idxUpdate_6[3:0]) begin
          TBEAddr_4 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEAddr_4 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h4 == idxAlloc[3:0]) begin
              TBEAddr_4 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_4 <= _GEN_2027;
            end
          end else if (_T_177) begin
            if (4'h4 == idxUpdate_4[3:0]) begin
              TBEAddr_4 <= 32'h0;
            end else begin
              TBEAddr_4 <= _GEN_2027;
            end
          end else begin
            TBEAddr_4 <= _GEN_2027;
          end
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEAddr_4 <= 32'h0;
          end else begin
            TBEAddr_4 <= _GEN_2541;
          end
        end else begin
          TBEAddr_4 <= _GEN_2541;
        end
      end else if (isAlloc_5) begin
        if (4'h4 == idxAlloc[3:0]) begin
          TBEAddr_4 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_4 <= _GEN_2541;
        end
      end else if (_T_199) begin
        if (4'h4 == idxUpdate_5[3:0]) begin
          TBEAddr_4 <= 32'h0;
        end else begin
          TBEAddr_4 <= _GEN_2541;
        end
      end else begin
        TBEAddr_4 <= _GEN_2541;
      end
    end else if (_T_243) begin
      if (4'h4 == idxUpdate_7[3:0]) begin
        TBEAddr_4 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h4 == idxAlloc[3:0]) begin
          TBEAddr_4 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h4 == idxAlloc[3:0]) begin
            TBEAddr_4 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_4 <= _GEN_2541;
          end
        end else if (_T_199) begin
          if (4'h4 == idxUpdate_5[3:0]) begin
            TBEAddr_4 <= 32'h0;
          end else begin
            TBEAddr_4 <= _GEN_2541;
          end
        end else begin
          TBEAddr_4 <= _GEN_2541;
        end
      end else if (_T_221) begin
        if (4'h4 == idxUpdate_6[3:0]) begin
          TBEAddr_4 <= 32'h0;
        end else begin
          TBEAddr_4 <= _GEN_3055;
        end
      end else begin
        TBEAddr_4 <= _GEN_3055;
      end
    end else if (isAlloc_6) begin
      if (4'h4 == idxAlloc[3:0]) begin
        TBEAddr_4 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_4 <= _GEN_3055;
      end
    end else if (_T_221) begin
      if (4'h4 == idxUpdate_6[3:0]) begin
        TBEAddr_4 <= 32'h0;
      end else begin
        TBEAddr_4 <= _GEN_3055;
      end
    end else begin
      TBEAddr_4 <= _GEN_3055;
    end
    if (reset) begin
      TBEAddr_5 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h5 == idxAlloc[3:0]) begin
        TBEAddr_5 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'h5 == idxAlloc[3:0]) begin
          TBEAddr_5 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEAddr_5 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEAddr_5 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEAddr_5 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEAddr_5 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEAddr_5 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEAddr_5 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEAddr_5 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEAddr_5 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEAddr_5 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEAddr_5 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEAddr_5 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'h5 == idxUpdate_0[3:0]) begin
                    TBEAddr_5 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEAddr_5 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEAddr_5 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h5 == idxAlloc[3:0]) begin
                      TBEAddr_5 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h5 == idxUpdate_0[3:0]) begin
                      TBEAddr_5 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEAddr_5 <= 32'h0;
                  end else begin
                    TBEAddr_5 <= _GEN_486;
                  end
                end else begin
                  TBEAddr_5 <= _GEN_486;
                end
              end else if (isAlloc_1) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEAddr_5 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_5 <= _GEN_486;
                end
              end else if (_T_111) begin
                if (4'h5 == idxUpdate_1[3:0]) begin
                  TBEAddr_5 <= 32'h0;
                end else begin
                  TBEAddr_5 <= _GEN_486;
                end
              end else begin
                TBEAddr_5 <= _GEN_486;
              end
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEAddr_5 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEAddr_5 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h5 == idxAlloc[3:0]) begin
                    TBEAddr_5 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_5 <= _GEN_486;
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUpdate_1[3:0]) begin
                    TBEAddr_5 <= 32'h0;
                  end else begin
                    TBEAddr_5 <= _GEN_486;
                  end
                end else begin
                  TBEAddr_5 <= _GEN_486;
                end
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEAddr_5 <= 32'h0;
                end else begin
                  TBEAddr_5 <= _GEN_1000;
                end
              end else begin
                TBEAddr_5 <= _GEN_1000;
              end
            end else if (isAlloc_2) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEAddr_5 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_5 <= _GEN_1000;
              end
            end else if (_T_133) begin
              if (4'h5 == idxUpdate_2[3:0]) begin
                TBEAddr_5 <= 32'h0;
              end else begin
                TBEAddr_5 <= _GEN_1000;
              end
            end else begin
              TBEAddr_5 <= _GEN_1000;
            end
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEAddr_5 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEAddr_5 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h5 == idxAlloc[3:0]) begin
                  TBEAddr_5 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_5 <= _GEN_1000;
                end
              end else if (_T_133) begin
                if (4'h5 == idxUpdate_2[3:0]) begin
                  TBEAddr_5 <= 32'h0;
                end else begin
                  TBEAddr_5 <= _GEN_1000;
                end
              end else begin
                TBEAddr_5 <= _GEN_1000;
              end
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEAddr_5 <= 32'h0;
              end else begin
                TBEAddr_5 <= _GEN_1514;
              end
            end else begin
              TBEAddr_5 <= _GEN_1514;
            end
          end else if (isAlloc_3) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEAddr_5 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_5 <= _GEN_1514;
            end
          end else if (_T_155) begin
            if (4'h5 == idxUpdate_3[3:0]) begin
              TBEAddr_5 <= 32'h0;
            end else begin
              TBEAddr_5 <= _GEN_1514;
            end
          end else begin
            TBEAddr_5 <= _GEN_1514;
          end
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEAddr_5 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEAddr_5 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h5 == idxAlloc[3:0]) begin
                TBEAddr_5 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_5 <= _GEN_1514;
              end
            end else if (_T_155) begin
              if (4'h5 == idxUpdate_3[3:0]) begin
                TBEAddr_5 <= 32'h0;
              end else begin
                TBEAddr_5 <= _GEN_1514;
              end
            end else begin
              TBEAddr_5 <= _GEN_1514;
            end
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEAddr_5 <= 32'h0;
            end else begin
              TBEAddr_5 <= _GEN_2028;
            end
          end else begin
            TBEAddr_5 <= _GEN_2028;
          end
        end else if (isAlloc_4) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEAddr_5 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_5 <= _GEN_2028;
          end
        end else if (_T_177) begin
          if (4'h5 == idxUpdate_4[3:0]) begin
            TBEAddr_5 <= 32'h0;
          end else begin
            TBEAddr_5 <= _GEN_2028;
          end
        end else begin
          TBEAddr_5 <= _GEN_2028;
        end
      end else if (_T_221) begin
        if (4'h5 == idxUpdate_6[3:0]) begin
          TBEAddr_5 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEAddr_5 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h5 == idxAlloc[3:0]) begin
              TBEAddr_5 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_5 <= _GEN_2028;
            end
          end else if (_T_177) begin
            if (4'h5 == idxUpdate_4[3:0]) begin
              TBEAddr_5 <= 32'h0;
            end else begin
              TBEAddr_5 <= _GEN_2028;
            end
          end else begin
            TBEAddr_5 <= _GEN_2028;
          end
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEAddr_5 <= 32'h0;
          end else begin
            TBEAddr_5 <= _GEN_2542;
          end
        end else begin
          TBEAddr_5 <= _GEN_2542;
        end
      end else if (isAlloc_5) begin
        if (4'h5 == idxAlloc[3:0]) begin
          TBEAddr_5 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_5 <= _GEN_2542;
        end
      end else if (_T_199) begin
        if (4'h5 == idxUpdate_5[3:0]) begin
          TBEAddr_5 <= 32'h0;
        end else begin
          TBEAddr_5 <= _GEN_2542;
        end
      end else begin
        TBEAddr_5 <= _GEN_2542;
      end
    end else if (_T_243) begin
      if (4'h5 == idxUpdate_7[3:0]) begin
        TBEAddr_5 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h5 == idxAlloc[3:0]) begin
          TBEAddr_5 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h5 == idxAlloc[3:0]) begin
            TBEAddr_5 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_5 <= _GEN_2542;
          end
        end else if (_T_199) begin
          if (4'h5 == idxUpdate_5[3:0]) begin
            TBEAddr_5 <= 32'h0;
          end else begin
            TBEAddr_5 <= _GEN_2542;
          end
        end else begin
          TBEAddr_5 <= _GEN_2542;
        end
      end else if (_T_221) begin
        if (4'h5 == idxUpdate_6[3:0]) begin
          TBEAddr_5 <= 32'h0;
        end else begin
          TBEAddr_5 <= _GEN_3056;
        end
      end else begin
        TBEAddr_5 <= _GEN_3056;
      end
    end else if (isAlloc_6) begin
      if (4'h5 == idxAlloc[3:0]) begin
        TBEAddr_5 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_5 <= _GEN_3056;
      end
    end else if (_T_221) begin
      if (4'h5 == idxUpdate_6[3:0]) begin
        TBEAddr_5 <= 32'h0;
      end else begin
        TBEAddr_5 <= _GEN_3056;
      end
    end else begin
      TBEAddr_5 <= _GEN_3056;
    end
    if (reset) begin
      TBEAddr_6 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h6 == idxAlloc[3:0]) begin
        TBEAddr_6 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'h6 == idxAlloc[3:0]) begin
          TBEAddr_6 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEAddr_6 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEAddr_6 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEAddr_6 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEAddr_6 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEAddr_6 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEAddr_6 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEAddr_6 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEAddr_6 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEAddr_6 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEAddr_6 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEAddr_6 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'h6 == idxUpdate_0[3:0]) begin
                    TBEAddr_6 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEAddr_6 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEAddr_6 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h6 == idxAlloc[3:0]) begin
                      TBEAddr_6 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h6 == idxUpdate_0[3:0]) begin
                      TBEAddr_6 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEAddr_6 <= 32'h0;
                  end else begin
                    TBEAddr_6 <= _GEN_487;
                  end
                end else begin
                  TBEAddr_6 <= _GEN_487;
                end
              end else if (isAlloc_1) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEAddr_6 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_6 <= _GEN_487;
                end
              end else if (_T_111) begin
                if (4'h6 == idxUpdate_1[3:0]) begin
                  TBEAddr_6 <= 32'h0;
                end else begin
                  TBEAddr_6 <= _GEN_487;
                end
              end else begin
                TBEAddr_6 <= _GEN_487;
              end
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEAddr_6 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEAddr_6 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h6 == idxAlloc[3:0]) begin
                    TBEAddr_6 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_6 <= _GEN_487;
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUpdate_1[3:0]) begin
                    TBEAddr_6 <= 32'h0;
                  end else begin
                    TBEAddr_6 <= _GEN_487;
                  end
                end else begin
                  TBEAddr_6 <= _GEN_487;
                end
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEAddr_6 <= 32'h0;
                end else begin
                  TBEAddr_6 <= _GEN_1001;
                end
              end else begin
                TBEAddr_6 <= _GEN_1001;
              end
            end else if (isAlloc_2) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEAddr_6 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_6 <= _GEN_1001;
              end
            end else if (_T_133) begin
              if (4'h6 == idxUpdate_2[3:0]) begin
                TBEAddr_6 <= 32'h0;
              end else begin
                TBEAddr_6 <= _GEN_1001;
              end
            end else begin
              TBEAddr_6 <= _GEN_1001;
            end
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEAddr_6 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEAddr_6 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h6 == idxAlloc[3:0]) begin
                  TBEAddr_6 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_6 <= _GEN_1001;
                end
              end else if (_T_133) begin
                if (4'h6 == idxUpdate_2[3:0]) begin
                  TBEAddr_6 <= 32'h0;
                end else begin
                  TBEAddr_6 <= _GEN_1001;
                end
              end else begin
                TBEAddr_6 <= _GEN_1001;
              end
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEAddr_6 <= 32'h0;
              end else begin
                TBEAddr_6 <= _GEN_1515;
              end
            end else begin
              TBEAddr_6 <= _GEN_1515;
            end
          end else if (isAlloc_3) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEAddr_6 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_6 <= _GEN_1515;
            end
          end else if (_T_155) begin
            if (4'h6 == idxUpdate_3[3:0]) begin
              TBEAddr_6 <= 32'h0;
            end else begin
              TBEAddr_6 <= _GEN_1515;
            end
          end else begin
            TBEAddr_6 <= _GEN_1515;
          end
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEAddr_6 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEAddr_6 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h6 == idxAlloc[3:0]) begin
                TBEAddr_6 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_6 <= _GEN_1515;
              end
            end else if (_T_155) begin
              if (4'h6 == idxUpdate_3[3:0]) begin
                TBEAddr_6 <= 32'h0;
              end else begin
                TBEAddr_6 <= _GEN_1515;
              end
            end else begin
              TBEAddr_6 <= _GEN_1515;
            end
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEAddr_6 <= 32'h0;
            end else begin
              TBEAddr_6 <= _GEN_2029;
            end
          end else begin
            TBEAddr_6 <= _GEN_2029;
          end
        end else if (isAlloc_4) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEAddr_6 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_6 <= _GEN_2029;
          end
        end else if (_T_177) begin
          if (4'h6 == idxUpdate_4[3:0]) begin
            TBEAddr_6 <= 32'h0;
          end else begin
            TBEAddr_6 <= _GEN_2029;
          end
        end else begin
          TBEAddr_6 <= _GEN_2029;
        end
      end else if (_T_221) begin
        if (4'h6 == idxUpdate_6[3:0]) begin
          TBEAddr_6 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEAddr_6 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h6 == idxAlloc[3:0]) begin
              TBEAddr_6 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_6 <= _GEN_2029;
            end
          end else if (_T_177) begin
            if (4'h6 == idxUpdate_4[3:0]) begin
              TBEAddr_6 <= 32'h0;
            end else begin
              TBEAddr_6 <= _GEN_2029;
            end
          end else begin
            TBEAddr_6 <= _GEN_2029;
          end
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEAddr_6 <= 32'h0;
          end else begin
            TBEAddr_6 <= _GEN_2543;
          end
        end else begin
          TBEAddr_6 <= _GEN_2543;
        end
      end else if (isAlloc_5) begin
        if (4'h6 == idxAlloc[3:0]) begin
          TBEAddr_6 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_6 <= _GEN_2543;
        end
      end else if (_T_199) begin
        if (4'h6 == idxUpdate_5[3:0]) begin
          TBEAddr_6 <= 32'h0;
        end else begin
          TBEAddr_6 <= _GEN_2543;
        end
      end else begin
        TBEAddr_6 <= _GEN_2543;
      end
    end else if (_T_243) begin
      if (4'h6 == idxUpdate_7[3:0]) begin
        TBEAddr_6 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h6 == idxAlloc[3:0]) begin
          TBEAddr_6 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h6 == idxAlloc[3:0]) begin
            TBEAddr_6 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_6 <= _GEN_2543;
          end
        end else if (_T_199) begin
          if (4'h6 == idxUpdate_5[3:0]) begin
            TBEAddr_6 <= 32'h0;
          end else begin
            TBEAddr_6 <= _GEN_2543;
          end
        end else begin
          TBEAddr_6 <= _GEN_2543;
        end
      end else if (_T_221) begin
        if (4'h6 == idxUpdate_6[3:0]) begin
          TBEAddr_6 <= 32'h0;
        end else begin
          TBEAddr_6 <= _GEN_3057;
        end
      end else begin
        TBEAddr_6 <= _GEN_3057;
      end
    end else if (isAlloc_6) begin
      if (4'h6 == idxAlloc[3:0]) begin
        TBEAddr_6 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_6 <= _GEN_3057;
      end
    end else if (_T_221) begin
      if (4'h6 == idxUpdate_6[3:0]) begin
        TBEAddr_6 <= 32'h0;
      end else begin
        TBEAddr_6 <= _GEN_3057;
      end
    end else begin
      TBEAddr_6 <= _GEN_3057;
    end
    if (reset) begin
      TBEAddr_7 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h7 == idxAlloc[3:0]) begin
        TBEAddr_7 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'h7 == idxAlloc[3:0]) begin
          TBEAddr_7 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEAddr_7 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEAddr_7 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEAddr_7 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEAddr_7 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEAddr_7 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEAddr_7 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEAddr_7 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEAddr_7 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEAddr_7 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEAddr_7 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEAddr_7 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'h7 == idxUpdate_0[3:0]) begin
                    TBEAddr_7 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEAddr_7 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEAddr_7 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h7 == idxAlloc[3:0]) begin
                      TBEAddr_7 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h7 == idxUpdate_0[3:0]) begin
                      TBEAddr_7 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEAddr_7 <= 32'h0;
                  end else begin
                    TBEAddr_7 <= _GEN_488;
                  end
                end else begin
                  TBEAddr_7 <= _GEN_488;
                end
              end else if (isAlloc_1) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEAddr_7 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_7 <= _GEN_488;
                end
              end else if (_T_111) begin
                if (4'h7 == idxUpdate_1[3:0]) begin
                  TBEAddr_7 <= 32'h0;
                end else begin
                  TBEAddr_7 <= _GEN_488;
                end
              end else begin
                TBEAddr_7 <= _GEN_488;
              end
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEAddr_7 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEAddr_7 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h7 == idxAlloc[3:0]) begin
                    TBEAddr_7 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_7 <= _GEN_488;
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUpdate_1[3:0]) begin
                    TBEAddr_7 <= 32'h0;
                  end else begin
                    TBEAddr_7 <= _GEN_488;
                  end
                end else begin
                  TBEAddr_7 <= _GEN_488;
                end
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEAddr_7 <= 32'h0;
                end else begin
                  TBEAddr_7 <= _GEN_1002;
                end
              end else begin
                TBEAddr_7 <= _GEN_1002;
              end
            end else if (isAlloc_2) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEAddr_7 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_7 <= _GEN_1002;
              end
            end else if (_T_133) begin
              if (4'h7 == idxUpdate_2[3:0]) begin
                TBEAddr_7 <= 32'h0;
              end else begin
                TBEAddr_7 <= _GEN_1002;
              end
            end else begin
              TBEAddr_7 <= _GEN_1002;
            end
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEAddr_7 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEAddr_7 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h7 == idxAlloc[3:0]) begin
                  TBEAddr_7 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_7 <= _GEN_1002;
                end
              end else if (_T_133) begin
                if (4'h7 == idxUpdate_2[3:0]) begin
                  TBEAddr_7 <= 32'h0;
                end else begin
                  TBEAddr_7 <= _GEN_1002;
                end
              end else begin
                TBEAddr_7 <= _GEN_1002;
              end
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEAddr_7 <= 32'h0;
              end else begin
                TBEAddr_7 <= _GEN_1516;
              end
            end else begin
              TBEAddr_7 <= _GEN_1516;
            end
          end else if (isAlloc_3) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEAddr_7 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_7 <= _GEN_1516;
            end
          end else if (_T_155) begin
            if (4'h7 == idxUpdate_3[3:0]) begin
              TBEAddr_7 <= 32'h0;
            end else begin
              TBEAddr_7 <= _GEN_1516;
            end
          end else begin
            TBEAddr_7 <= _GEN_1516;
          end
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEAddr_7 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEAddr_7 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h7 == idxAlloc[3:0]) begin
                TBEAddr_7 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_7 <= _GEN_1516;
              end
            end else if (_T_155) begin
              if (4'h7 == idxUpdate_3[3:0]) begin
                TBEAddr_7 <= 32'h0;
              end else begin
                TBEAddr_7 <= _GEN_1516;
              end
            end else begin
              TBEAddr_7 <= _GEN_1516;
            end
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEAddr_7 <= 32'h0;
            end else begin
              TBEAddr_7 <= _GEN_2030;
            end
          end else begin
            TBEAddr_7 <= _GEN_2030;
          end
        end else if (isAlloc_4) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEAddr_7 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_7 <= _GEN_2030;
          end
        end else if (_T_177) begin
          if (4'h7 == idxUpdate_4[3:0]) begin
            TBEAddr_7 <= 32'h0;
          end else begin
            TBEAddr_7 <= _GEN_2030;
          end
        end else begin
          TBEAddr_7 <= _GEN_2030;
        end
      end else if (_T_221) begin
        if (4'h7 == idxUpdate_6[3:0]) begin
          TBEAddr_7 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEAddr_7 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h7 == idxAlloc[3:0]) begin
              TBEAddr_7 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_7 <= _GEN_2030;
            end
          end else if (_T_177) begin
            if (4'h7 == idxUpdate_4[3:0]) begin
              TBEAddr_7 <= 32'h0;
            end else begin
              TBEAddr_7 <= _GEN_2030;
            end
          end else begin
            TBEAddr_7 <= _GEN_2030;
          end
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEAddr_7 <= 32'h0;
          end else begin
            TBEAddr_7 <= _GEN_2544;
          end
        end else begin
          TBEAddr_7 <= _GEN_2544;
        end
      end else if (isAlloc_5) begin
        if (4'h7 == idxAlloc[3:0]) begin
          TBEAddr_7 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_7 <= _GEN_2544;
        end
      end else if (_T_199) begin
        if (4'h7 == idxUpdate_5[3:0]) begin
          TBEAddr_7 <= 32'h0;
        end else begin
          TBEAddr_7 <= _GEN_2544;
        end
      end else begin
        TBEAddr_7 <= _GEN_2544;
      end
    end else if (_T_243) begin
      if (4'h7 == idxUpdate_7[3:0]) begin
        TBEAddr_7 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h7 == idxAlloc[3:0]) begin
          TBEAddr_7 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h7 == idxAlloc[3:0]) begin
            TBEAddr_7 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_7 <= _GEN_2544;
          end
        end else if (_T_199) begin
          if (4'h7 == idxUpdate_5[3:0]) begin
            TBEAddr_7 <= 32'h0;
          end else begin
            TBEAddr_7 <= _GEN_2544;
          end
        end else begin
          TBEAddr_7 <= _GEN_2544;
        end
      end else if (_T_221) begin
        if (4'h7 == idxUpdate_6[3:0]) begin
          TBEAddr_7 <= 32'h0;
        end else begin
          TBEAddr_7 <= _GEN_3058;
        end
      end else begin
        TBEAddr_7 <= _GEN_3058;
      end
    end else if (isAlloc_6) begin
      if (4'h7 == idxAlloc[3:0]) begin
        TBEAddr_7 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_7 <= _GEN_3058;
      end
    end else if (_T_221) begin
      if (4'h7 == idxUpdate_6[3:0]) begin
        TBEAddr_7 <= 32'h0;
      end else begin
        TBEAddr_7 <= _GEN_3058;
      end
    end else begin
      TBEAddr_7 <= _GEN_3058;
    end
    if (reset) begin
      TBEAddr_8 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h8 == idxAlloc[3:0]) begin
        TBEAddr_8 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'h8 == idxAlloc[3:0]) begin
          TBEAddr_8 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEAddr_8 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEAddr_8 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEAddr_8 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEAddr_8 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEAddr_8 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEAddr_8 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEAddr_8 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEAddr_8 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEAddr_8 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEAddr_8 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEAddr_8 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'h8 == idxUpdate_0[3:0]) begin
                    TBEAddr_8 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEAddr_8 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEAddr_8 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h8 == idxAlloc[3:0]) begin
                      TBEAddr_8 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h8 == idxUpdate_0[3:0]) begin
                      TBEAddr_8 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEAddr_8 <= 32'h0;
                  end else begin
                    TBEAddr_8 <= _GEN_489;
                  end
                end else begin
                  TBEAddr_8 <= _GEN_489;
                end
              end else if (isAlloc_1) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEAddr_8 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_8 <= _GEN_489;
                end
              end else if (_T_111) begin
                if (4'h8 == idxUpdate_1[3:0]) begin
                  TBEAddr_8 <= 32'h0;
                end else begin
                  TBEAddr_8 <= _GEN_489;
                end
              end else begin
                TBEAddr_8 <= _GEN_489;
              end
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEAddr_8 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEAddr_8 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h8 == idxAlloc[3:0]) begin
                    TBEAddr_8 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_8 <= _GEN_489;
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUpdate_1[3:0]) begin
                    TBEAddr_8 <= 32'h0;
                  end else begin
                    TBEAddr_8 <= _GEN_489;
                  end
                end else begin
                  TBEAddr_8 <= _GEN_489;
                end
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEAddr_8 <= 32'h0;
                end else begin
                  TBEAddr_8 <= _GEN_1003;
                end
              end else begin
                TBEAddr_8 <= _GEN_1003;
              end
            end else if (isAlloc_2) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEAddr_8 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_8 <= _GEN_1003;
              end
            end else if (_T_133) begin
              if (4'h8 == idxUpdate_2[3:0]) begin
                TBEAddr_8 <= 32'h0;
              end else begin
                TBEAddr_8 <= _GEN_1003;
              end
            end else begin
              TBEAddr_8 <= _GEN_1003;
            end
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEAddr_8 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEAddr_8 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h8 == idxAlloc[3:0]) begin
                  TBEAddr_8 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_8 <= _GEN_1003;
                end
              end else if (_T_133) begin
                if (4'h8 == idxUpdate_2[3:0]) begin
                  TBEAddr_8 <= 32'h0;
                end else begin
                  TBEAddr_8 <= _GEN_1003;
                end
              end else begin
                TBEAddr_8 <= _GEN_1003;
              end
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEAddr_8 <= 32'h0;
              end else begin
                TBEAddr_8 <= _GEN_1517;
              end
            end else begin
              TBEAddr_8 <= _GEN_1517;
            end
          end else if (isAlloc_3) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEAddr_8 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_8 <= _GEN_1517;
            end
          end else if (_T_155) begin
            if (4'h8 == idxUpdate_3[3:0]) begin
              TBEAddr_8 <= 32'h0;
            end else begin
              TBEAddr_8 <= _GEN_1517;
            end
          end else begin
            TBEAddr_8 <= _GEN_1517;
          end
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEAddr_8 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEAddr_8 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h8 == idxAlloc[3:0]) begin
                TBEAddr_8 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_8 <= _GEN_1517;
              end
            end else if (_T_155) begin
              if (4'h8 == idxUpdate_3[3:0]) begin
                TBEAddr_8 <= 32'h0;
              end else begin
                TBEAddr_8 <= _GEN_1517;
              end
            end else begin
              TBEAddr_8 <= _GEN_1517;
            end
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEAddr_8 <= 32'h0;
            end else begin
              TBEAddr_8 <= _GEN_2031;
            end
          end else begin
            TBEAddr_8 <= _GEN_2031;
          end
        end else if (isAlloc_4) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEAddr_8 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_8 <= _GEN_2031;
          end
        end else if (_T_177) begin
          if (4'h8 == idxUpdate_4[3:0]) begin
            TBEAddr_8 <= 32'h0;
          end else begin
            TBEAddr_8 <= _GEN_2031;
          end
        end else begin
          TBEAddr_8 <= _GEN_2031;
        end
      end else if (_T_221) begin
        if (4'h8 == idxUpdate_6[3:0]) begin
          TBEAddr_8 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEAddr_8 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h8 == idxAlloc[3:0]) begin
              TBEAddr_8 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_8 <= _GEN_2031;
            end
          end else if (_T_177) begin
            if (4'h8 == idxUpdate_4[3:0]) begin
              TBEAddr_8 <= 32'h0;
            end else begin
              TBEAddr_8 <= _GEN_2031;
            end
          end else begin
            TBEAddr_8 <= _GEN_2031;
          end
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEAddr_8 <= 32'h0;
          end else begin
            TBEAddr_8 <= _GEN_2545;
          end
        end else begin
          TBEAddr_8 <= _GEN_2545;
        end
      end else if (isAlloc_5) begin
        if (4'h8 == idxAlloc[3:0]) begin
          TBEAddr_8 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_8 <= _GEN_2545;
        end
      end else if (_T_199) begin
        if (4'h8 == idxUpdate_5[3:0]) begin
          TBEAddr_8 <= 32'h0;
        end else begin
          TBEAddr_8 <= _GEN_2545;
        end
      end else begin
        TBEAddr_8 <= _GEN_2545;
      end
    end else if (_T_243) begin
      if (4'h8 == idxUpdate_7[3:0]) begin
        TBEAddr_8 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h8 == idxAlloc[3:0]) begin
          TBEAddr_8 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h8 == idxAlloc[3:0]) begin
            TBEAddr_8 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_8 <= _GEN_2545;
          end
        end else if (_T_199) begin
          if (4'h8 == idxUpdate_5[3:0]) begin
            TBEAddr_8 <= 32'h0;
          end else begin
            TBEAddr_8 <= _GEN_2545;
          end
        end else begin
          TBEAddr_8 <= _GEN_2545;
        end
      end else if (_T_221) begin
        if (4'h8 == idxUpdate_6[3:0]) begin
          TBEAddr_8 <= 32'h0;
        end else begin
          TBEAddr_8 <= _GEN_3059;
        end
      end else begin
        TBEAddr_8 <= _GEN_3059;
      end
    end else if (isAlloc_6) begin
      if (4'h8 == idxAlloc[3:0]) begin
        TBEAddr_8 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_8 <= _GEN_3059;
      end
    end else if (_T_221) begin
      if (4'h8 == idxUpdate_6[3:0]) begin
        TBEAddr_8 <= 32'h0;
      end else begin
        TBEAddr_8 <= _GEN_3059;
      end
    end else begin
      TBEAddr_8 <= _GEN_3059;
    end
    if (reset) begin
      TBEAddr_9 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'h9 == idxAlloc[3:0]) begin
        TBEAddr_9 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'h9 == idxAlloc[3:0]) begin
          TBEAddr_9 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEAddr_9 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEAddr_9 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEAddr_9 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEAddr_9 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEAddr_9 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEAddr_9 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEAddr_9 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEAddr_9 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEAddr_9 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEAddr_9 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEAddr_9 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'h9 == idxUpdate_0[3:0]) begin
                    TBEAddr_9 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEAddr_9 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEAddr_9 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'h9 == idxAlloc[3:0]) begin
                      TBEAddr_9 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'h9 == idxUpdate_0[3:0]) begin
                      TBEAddr_9 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEAddr_9 <= 32'h0;
                  end else begin
                    TBEAddr_9 <= _GEN_490;
                  end
                end else begin
                  TBEAddr_9 <= _GEN_490;
                end
              end else if (isAlloc_1) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEAddr_9 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_9 <= _GEN_490;
                end
              end else if (_T_111) begin
                if (4'h9 == idxUpdate_1[3:0]) begin
                  TBEAddr_9 <= 32'h0;
                end else begin
                  TBEAddr_9 <= _GEN_490;
                end
              end else begin
                TBEAddr_9 <= _GEN_490;
              end
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEAddr_9 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEAddr_9 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'h9 == idxAlloc[3:0]) begin
                    TBEAddr_9 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_9 <= _GEN_490;
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUpdate_1[3:0]) begin
                    TBEAddr_9 <= 32'h0;
                  end else begin
                    TBEAddr_9 <= _GEN_490;
                  end
                end else begin
                  TBEAddr_9 <= _GEN_490;
                end
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEAddr_9 <= 32'h0;
                end else begin
                  TBEAddr_9 <= _GEN_1004;
                end
              end else begin
                TBEAddr_9 <= _GEN_1004;
              end
            end else if (isAlloc_2) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEAddr_9 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_9 <= _GEN_1004;
              end
            end else if (_T_133) begin
              if (4'h9 == idxUpdate_2[3:0]) begin
                TBEAddr_9 <= 32'h0;
              end else begin
                TBEAddr_9 <= _GEN_1004;
              end
            end else begin
              TBEAddr_9 <= _GEN_1004;
            end
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEAddr_9 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEAddr_9 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'h9 == idxAlloc[3:0]) begin
                  TBEAddr_9 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_9 <= _GEN_1004;
                end
              end else if (_T_133) begin
                if (4'h9 == idxUpdate_2[3:0]) begin
                  TBEAddr_9 <= 32'h0;
                end else begin
                  TBEAddr_9 <= _GEN_1004;
                end
              end else begin
                TBEAddr_9 <= _GEN_1004;
              end
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEAddr_9 <= 32'h0;
              end else begin
                TBEAddr_9 <= _GEN_1518;
              end
            end else begin
              TBEAddr_9 <= _GEN_1518;
            end
          end else if (isAlloc_3) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEAddr_9 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_9 <= _GEN_1518;
            end
          end else if (_T_155) begin
            if (4'h9 == idxUpdate_3[3:0]) begin
              TBEAddr_9 <= 32'h0;
            end else begin
              TBEAddr_9 <= _GEN_1518;
            end
          end else begin
            TBEAddr_9 <= _GEN_1518;
          end
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEAddr_9 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEAddr_9 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'h9 == idxAlloc[3:0]) begin
                TBEAddr_9 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_9 <= _GEN_1518;
              end
            end else if (_T_155) begin
              if (4'h9 == idxUpdate_3[3:0]) begin
                TBEAddr_9 <= 32'h0;
              end else begin
                TBEAddr_9 <= _GEN_1518;
              end
            end else begin
              TBEAddr_9 <= _GEN_1518;
            end
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEAddr_9 <= 32'h0;
            end else begin
              TBEAddr_9 <= _GEN_2032;
            end
          end else begin
            TBEAddr_9 <= _GEN_2032;
          end
        end else if (isAlloc_4) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEAddr_9 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_9 <= _GEN_2032;
          end
        end else if (_T_177) begin
          if (4'h9 == idxUpdate_4[3:0]) begin
            TBEAddr_9 <= 32'h0;
          end else begin
            TBEAddr_9 <= _GEN_2032;
          end
        end else begin
          TBEAddr_9 <= _GEN_2032;
        end
      end else if (_T_221) begin
        if (4'h9 == idxUpdate_6[3:0]) begin
          TBEAddr_9 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEAddr_9 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'h9 == idxAlloc[3:0]) begin
              TBEAddr_9 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_9 <= _GEN_2032;
            end
          end else if (_T_177) begin
            if (4'h9 == idxUpdate_4[3:0]) begin
              TBEAddr_9 <= 32'h0;
            end else begin
              TBEAddr_9 <= _GEN_2032;
            end
          end else begin
            TBEAddr_9 <= _GEN_2032;
          end
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEAddr_9 <= 32'h0;
          end else begin
            TBEAddr_9 <= _GEN_2546;
          end
        end else begin
          TBEAddr_9 <= _GEN_2546;
        end
      end else if (isAlloc_5) begin
        if (4'h9 == idxAlloc[3:0]) begin
          TBEAddr_9 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_9 <= _GEN_2546;
        end
      end else if (_T_199) begin
        if (4'h9 == idxUpdate_5[3:0]) begin
          TBEAddr_9 <= 32'h0;
        end else begin
          TBEAddr_9 <= _GEN_2546;
        end
      end else begin
        TBEAddr_9 <= _GEN_2546;
      end
    end else if (_T_243) begin
      if (4'h9 == idxUpdate_7[3:0]) begin
        TBEAddr_9 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'h9 == idxAlloc[3:0]) begin
          TBEAddr_9 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'h9 == idxAlloc[3:0]) begin
            TBEAddr_9 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_9 <= _GEN_2546;
          end
        end else if (_T_199) begin
          if (4'h9 == idxUpdate_5[3:0]) begin
            TBEAddr_9 <= 32'h0;
          end else begin
            TBEAddr_9 <= _GEN_2546;
          end
        end else begin
          TBEAddr_9 <= _GEN_2546;
        end
      end else if (_T_221) begin
        if (4'h9 == idxUpdate_6[3:0]) begin
          TBEAddr_9 <= 32'h0;
        end else begin
          TBEAddr_9 <= _GEN_3060;
        end
      end else begin
        TBEAddr_9 <= _GEN_3060;
      end
    end else if (isAlloc_6) begin
      if (4'h9 == idxAlloc[3:0]) begin
        TBEAddr_9 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_9 <= _GEN_3060;
      end
    end else if (_T_221) begin
      if (4'h9 == idxUpdate_6[3:0]) begin
        TBEAddr_9 <= 32'h0;
      end else begin
        TBEAddr_9 <= _GEN_3060;
      end
    end else begin
      TBEAddr_9 <= _GEN_3060;
    end
    if (reset) begin
      TBEAddr_10 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'ha == idxAlloc[3:0]) begin
        TBEAddr_10 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'ha == idxAlloc[3:0]) begin
          TBEAddr_10 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEAddr_10 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEAddr_10 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEAddr_10 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEAddr_10 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEAddr_10 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEAddr_10 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEAddr_10 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEAddr_10 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEAddr_10 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEAddr_10 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEAddr_10 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'ha == idxUpdate_0[3:0]) begin
                    TBEAddr_10 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEAddr_10 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEAddr_10 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'ha == idxAlloc[3:0]) begin
                      TBEAddr_10 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'ha == idxUpdate_0[3:0]) begin
                      TBEAddr_10 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEAddr_10 <= 32'h0;
                  end else begin
                    TBEAddr_10 <= _GEN_491;
                  end
                end else begin
                  TBEAddr_10 <= _GEN_491;
                end
              end else if (isAlloc_1) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEAddr_10 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_10 <= _GEN_491;
                end
              end else if (_T_111) begin
                if (4'ha == idxUpdate_1[3:0]) begin
                  TBEAddr_10 <= 32'h0;
                end else begin
                  TBEAddr_10 <= _GEN_491;
                end
              end else begin
                TBEAddr_10 <= _GEN_491;
              end
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEAddr_10 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEAddr_10 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'ha == idxAlloc[3:0]) begin
                    TBEAddr_10 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_10 <= _GEN_491;
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUpdate_1[3:0]) begin
                    TBEAddr_10 <= 32'h0;
                  end else begin
                    TBEAddr_10 <= _GEN_491;
                  end
                end else begin
                  TBEAddr_10 <= _GEN_491;
                end
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEAddr_10 <= 32'h0;
                end else begin
                  TBEAddr_10 <= _GEN_1005;
                end
              end else begin
                TBEAddr_10 <= _GEN_1005;
              end
            end else if (isAlloc_2) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEAddr_10 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_10 <= _GEN_1005;
              end
            end else if (_T_133) begin
              if (4'ha == idxUpdate_2[3:0]) begin
                TBEAddr_10 <= 32'h0;
              end else begin
                TBEAddr_10 <= _GEN_1005;
              end
            end else begin
              TBEAddr_10 <= _GEN_1005;
            end
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEAddr_10 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEAddr_10 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'ha == idxAlloc[3:0]) begin
                  TBEAddr_10 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_10 <= _GEN_1005;
                end
              end else if (_T_133) begin
                if (4'ha == idxUpdate_2[3:0]) begin
                  TBEAddr_10 <= 32'h0;
                end else begin
                  TBEAddr_10 <= _GEN_1005;
                end
              end else begin
                TBEAddr_10 <= _GEN_1005;
              end
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEAddr_10 <= 32'h0;
              end else begin
                TBEAddr_10 <= _GEN_1519;
              end
            end else begin
              TBEAddr_10 <= _GEN_1519;
            end
          end else if (isAlloc_3) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEAddr_10 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_10 <= _GEN_1519;
            end
          end else if (_T_155) begin
            if (4'ha == idxUpdate_3[3:0]) begin
              TBEAddr_10 <= 32'h0;
            end else begin
              TBEAddr_10 <= _GEN_1519;
            end
          end else begin
            TBEAddr_10 <= _GEN_1519;
          end
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEAddr_10 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEAddr_10 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'ha == idxAlloc[3:0]) begin
                TBEAddr_10 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_10 <= _GEN_1519;
              end
            end else if (_T_155) begin
              if (4'ha == idxUpdate_3[3:0]) begin
                TBEAddr_10 <= 32'h0;
              end else begin
                TBEAddr_10 <= _GEN_1519;
              end
            end else begin
              TBEAddr_10 <= _GEN_1519;
            end
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEAddr_10 <= 32'h0;
            end else begin
              TBEAddr_10 <= _GEN_2033;
            end
          end else begin
            TBEAddr_10 <= _GEN_2033;
          end
        end else if (isAlloc_4) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEAddr_10 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_10 <= _GEN_2033;
          end
        end else if (_T_177) begin
          if (4'ha == idxUpdate_4[3:0]) begin
            TBEAddr_10 <= 32'h0;
          end else begin
            TBEAddr_10 <= _GEN_2033;
          end
        end else begin
          TBEAddr_10 <= _GEN_2033;
        end
      end else if (_T_221) begin
        if (4'ha == idxUpdate_6[3:0]) begin
          TBEAddr_10 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEAddr_10 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'ha == idxAlloc[3:0]) begin
              TBEAddr_10 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_10 <= _GEN_2033;
            end
          end else if (_T_177) begin
            if (4'ha == idxUpdate_4[3:0]) begin
              TBEAddr_10 <= 32'h0;
            end else begin
              TBEAddr_10 <= _GEN_2033;
            end
          end else begin
            TBEAddr_10 <= _GEN_2033;
          end
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEAddr_10 <= 32'h0;
          end else begin
            TBEAddr_10 <= _GEN_2547;
          end
        end else begin
          TBEAddr_10 <= _GEN_2547;
        end
      end else if (isAlloc_5) begin
        if (4'ha == idxAlloc[3:0]) begin
          TBEAddr_10 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_10 <= _GEN_2547;
        end
      end else if (_T_199) begin
        if (4'ha == idxUpdate_5[3:0]) begin
          TBEAddr_10 <= 32'h0;
        end else begin
          TBEAddr_10 <= _GEN_2547;
        end
      end else begin
        TBEAddr_10 <= _GEN_2547;
      end
    end else if (_T_243) begin
      if (4'ha == idxUpdate_7[3:0]) begin
        TBEAddr_10 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'ha == idxAlloc[3:0]) begin
          TBEAddr_10 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'ha == idxAlloc[3:0]) begin
            TBEAddr_10 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_10 <= _GEN_2547;
          end
        end else if (_T_199) begin
          if (4'ha == idxUpdate_5[3:0]) begin
            TBEAddr_10 <= 32'h0;
          end else begin
            TBEAddr_10 <= _GEN_2547;
          end
        end else begin
          TBEAddr_10 <= _GEN_2547;
        end
      end else if (_T_221) begin
        if (4'ha == idxUpdate_6[3:0]) begin
          TBEAddr_10 <= 32'h0;
        end else begin
          TBEAddr_10 <= _GEN_3061;
        end
      end else begin
        TBEAddr_10 <= _GEN_3061;
      end
    end else if (isAlloc_6) begin
      if (4'ha == idxAlloc[3:0]) begin
        TBEAddr_10 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_10 <= _GEN_3061;
      end
    end else if (_T_221) begin
      if (4'ha == idxUpdate_6[3:0]) begin
        TBEAddr_10 <= 32'h0;
      end else begin
        TBEAddr_10 <= _GEN_3061;
      end
    end else begin
      TBEAddr_10 <= _GEN_3061;
    end
    if (reset) begin
      TBEAddr_11 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'hb == idxAlloc[3:0]) begin
        TBEAddr_11 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'hb == idxAlloc[3:0]) begin
          TBEAddr_11 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEAddr_11 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEAddr_11 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEAddr_11 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEAddr_11 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEAddr_11 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEAddr_11 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEAddr_11 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEAddr_11 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEAddr_11 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEAddr_11 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEAddr_11 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'hb == idxUpdate_0[3:0]) begin
                    TBEAddr_11 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEAddr_11 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEAddr_11 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'hb == idxAlloc[3:0]) begin
                      TBEAddr_11 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'hb == idxUpdate_0[3:0]) begin
                      TBEAddr_11 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEAddr_11 <= 32'h0;
                  end else begin
                    TBEAddr_11 <= _GEN_492;
                  end
                end else begin
                  TBEAddr_11 <= _GEN_492;
                end
              end else if (isAlloc_1) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEAddr_11 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_11 <= _GEN_492;
                end
              end else if (_T_111) begin
                if (4'hb == idxUpdate_1[3:0]) begin
                  TBEAddr_11 <= 32'h0;
                end else begin
                  TBEAddr_11 <= _GEN_492;
                end
              end else begin
                TBEAddr_11 <= _GEN_492;
              end
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEAddr_11 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEAddr_11 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'hb == idxAlloc[3:0]) begin
                    TBEAddr_11 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_11 <= _GEN_492;
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUpdate_1[3:0]) begin
                    TBEAddr_11 <= 32'h0;
                  end else begin
                    TBEAddr_11 <= _GEN_492;
                  end
                end else begin
                  TBEAddr_11 <= _GEN_492;
                end
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEAddr_11 <= 32'h0;
                end else begin
                  TBEAddr_11 <= _GEN_1006;
                end
              end else begin
                TBEAddr_11 <= _GEN_1006;
              end
            end else if (isAlloc_2) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEAddr_11 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_11 <= _GEN_1006;
              end
            end else if (_T_133) begin
              if (4'hb == idxUpdate_2[3:0]) begin
                TBEAddr_11 <= 32'h0;
              end else begin
                TBEAddr_11 <= _GEN_1006;
              end
            end else begin
              TBEAddr_11 <= _GEN_1006;
            end
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEAddr_11 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEAddr_11 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'hb == idxAlloc[3:0]) begin
                  TBEAddr_11 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_11 <= _GEN_1006;
                end
              end else if (_T_133) begin
                if (4'hb == idxUpdate_2[3:0]) begin
                  TBEAddr_11 <= 32'h0;
                end else begin
                  TBEAddr_11 <= _GEN_1006;
                end
              end else begin
                TBEAddr_11 <= _GEN_1006;
              end
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEAddr_11 <= 32'h0;
              end else begin
                TBEAddr_11 <= _GEN_1520;
              end
            end else begin
              TBEAddr_11 <= _GEN_1520;
            end
          end else if (isAlloc_3) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEAddr_11 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_11 <= _GEN_1520;
            end
          end else if (_T_155) begin
            if (4'hb == idxUpdate_3[3:0]) begin
              TBEAddr_11 <= 32'h0;
            end else begin
              TBEAddr_11 <= _GEN_1520;
            end
          end else begin
            TBEAddr_11 <= _GEN_1520;
          end
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEAddr_11 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEAddr_11 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'hb == idxAlloc[3:0]) begin
                TBEAddr_11 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_11 <= _GEN_1520;
              end
            end else if (_T_155) begin
              if (4'hb == idxUpdate_3[3:0]) begin
                TBEAddr_11 <= 32'h0;
              end else begin
                TBEAddr_11 <= _GEN_1520;
              end
            end else begin
              TBEAddr_11 <= _GEN_1520;
            end
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEAddr_11 <= 32'h0;
            end else begin
              TBEAddr_11 <= _GEN_2034;
            end
          end else begin
            TBEAddr_11 <= _GEN_2034;
          end
        end else if (isAlloc_4) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEAddr_11 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_11 <= _GEN_2034;
          end
        end else if (_T_177) begin
          if (4'hb == idxUpdate_4[3:0]) begin
            TBEAddr_11 <= 32'h0;
          end else begin
            TBEAddr_11 <= _GEN_2034;
          end
        end else begin
          TBEAddr_11 <= _GEN_2034;
        end
      end else if (_T_221) begin
        if (4'hb == idxUpdate_6[3:0]) begin
          TBEAddr_11 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEAddr_11 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'hb == idxAlloc[3:0]) begin
              TBEAddr_11 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_11 <= _GEN_2034;
            end
          end else if (_T_177) begin
            if (4'hb == idxUpdate_4[3:0]) begin
              TBEAddr_11 <= 32'h0;
            end else begin
              TBEAddr_11 <= _GEN_2034;
            end
          end else begin
            TBEAddr_11 <= _GEN_2034;
          end
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEAddr_11 <= 32'h0;
          end else begin
            TBEAddr_11 <= _GEN_2548;
          end
        end else begin
          TBEAddr_11 <= _GEN_2548;
        end
      end else if (isAlloc_5) begin
        if (4'hb == idxAlloc[3:0]) begin
          TBEAddr_11 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_11 <= _GEN_2548;
        end
      end else if (_T_199) begin
        if (4'hb == idxUpdate_5[3:0]) begin
          TBEAddr_11 <= 32'h0;
        end else begin
          TBEAddr_11 <= _GEN_2548;
        end
      end else begin
        TBEAddr_11 <= _GEN_2548;
      end
    end else if (_T_243) begin
      if (4'hb == idxUpdate_7[3:0]) begin
        TBEAddr_11 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'hb == idxAlloc[3:0]) begin
          TBEAddr_11 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'hb == idxAlloc[3:0]) begin
            TBEAddr_11 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_11 <= _GEN_2548;
          end
        end else if (_T_199) begin
          if (4'hb == idxUpdate_5[3:0]) begin
            TBEAddr_11 <= 32'h0;
          end else begin
            TBEAddr_11 <= _GEN_2548;
          end
        end else begin
          TBEAddr_11 <= _GEN_2548;
        end
      end else if (_T_221) begin
        if (4'hb == idxUpdate_6[3:0]) begin
          TBEAddr_11 <= 32'h0;
        end else begin
          TBEAddr_11 <= _GEN_3062;
        end
      end else begin
        TBEAddr_11 <= _GEN_3062;
      end
    end else if (isAlloc_6) begin
      if (4'hb == idxAlloc[3:0]) begin
        TBEAddr_11 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_11 <= _GEN_3062;
      end
    end else if (_T_221) begin
      if (4'hb == idxUpdate_6[3:0]) begin
        TBEAddr_11 <= 32'h0;
      end else begin
        TBEAddr_11 <= _GEN_3062;
      end
    end else begin
      TBEAddr_11 <= _GEN_3062;
    end
    if (reset) begin
      TBEAddr_12 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'hc == idxAlloc[3:0]) begin
        TBEAddr_12 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'hc == idxAlloc[3:0]) begin
          TBEAddr_12 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEAddr_12 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEAddr_12 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEAddr_12 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEAddr_12 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEAddr_12 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEAddr_12 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEAddr_12 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEAddr_12 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEAddr_12 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEAddr_12 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEAddr_12 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'hc == idxUpdate_0[3:0]) begin
                    TBEAddr_12 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEAddr_12 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEAddr_12 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'hc == idxAlloc[3:0]) begin
                      TBEAddr_12 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'hc == idxUpdate_0[3:0]) begin
                      TBEAddr_12 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEAddr_12 <= 32'h0;
                  end else begin
                    TBEAddr_12 <= _GEN_493;
                  end
                end else begin
                  TBEAddr_12 <= _GEN_493;
                end
              end else if (isAlloc_1) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEAddr_12 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_12 <= _GEN_493;
                end
              end else if (_T_111) begin
                if (4'hc == idxUpdate_1[3:0]) begin
                  TBEAddr_12 <= 32'h0;
                end else begin
                  TBEAddr_12 <= _GEN_493;
                end
              end else begin
                TBEAddr_12 <= _GEN_493;
              end
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEAddr_12 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEAddr_12 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'hc == idxAlloc[3:0]) begin
                    TBEAddr_12 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_12 <= _GEN_493;
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUpdate_1[3:0]) begin
                    TBEAddr_12 <= 32'h0;
                  end else begin
                    TBEAddr_12 <= _GEN_493;
                  end
                end else begin
                  TBEAddr_12 <= _GEN_493;
                end
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEAddr_12 <= 32'h0;
                end else begin
                  TBEAddr_12 <= _GEN_1007;
                end
              end else begin
                TBEAddr_12 <= _GEN_1007;
              end
            end else if (isAlloc_2) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEAddr_12 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_12 <= _GEN_1007;
              end
            end else if (_T_133) begin
              if (4'hc == idxUpdate_2[3:0]) begin
                TBEAddr_12 <= 32'h0;
              end else begin
                TBEAddr_12 <= _GEN_1007;
              end
            end else begin
              TBEAddr_12 <= _GEN_1007;
            end
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEAddr_12 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEAddr_12 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'hc == idxAlloc[3:0]) begin
                  TBEAddr_12 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_12 <= _GEN_1007;
                end
              end else if (_T_133) begin
                if (4'hc == idxUpdate_2[3:0]) begin
                  TBEAddr_12 <= 32'h0;
                end else begin
                  TBEAddr_12 <= _GEN_1007;
                end
              end else begin
                TBEAddr_12 <= _GEN_1007;
              end
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEAddr_12 <= 32'h0;
              end else begin
                TBEAddr_12 <= _GEN_1521;
              end
            end else begin
              TBEAddr_12 <= _GEN_1521;
            end
          end else if (isAlloc_3) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEAddr_12 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_12 <= _GEN_1521;
            end
          end else if (_T_155) begin
            if (4'hc == idxUpdate_3[3:0]) begin
              TBEAddr_12 <= 32'h0;
            end else begin
              TBEAddr_12 <= _GEN_1521;
            end
          end else begin
            TBEAddr_12 <= _GEN_1521;
          end
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEAddr_12 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEAddr_12 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'hc == idxAlloc[3:0]) begin
                TBEAddr_12 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_12 <= _GEN_1521;
              end
            end else if (_T_155) begin
              if (4'hc == idxUpdate_3[3:0]) begin
                TBEAddr_12 <= 32'h0;
              end else begin
                TBEAddr_12 <= _GEN_1521;
              end
            end else begin
              TBEAddr_12 <= _GEN_1521;
            end
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEAddr_12 <= 32'h0;
            end else begin
              TBEAddr_12 <= _GEN_2035;
            end
          end else begin
            TBEAddr_12 <= _GEN_2035;
          end
        end else if (isAlloc_4) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEAddr_12 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_12 <= _GEN_2035;
          end
        end else if (_T_177) begin
          if (4'hc == idxUpdate_4[3:0]) begin
            TBEAddr_12 <= 32'h0;
          end else begin
            TBEAddr_12 <= _GEN_2035;
          end
        end else begin
          TBEAddr_12 <= _GEN_2035;
        end
      end else if (_T_221) begin
        if (4'hc == idxUpdate_6[3:0]) begin
          TBEAddr_12 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEAddr_12 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'hc == idxAlloc[3:0]) begin
              TBEAddr_12 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_12 <= _GEN_2035;
            end
          end else if (_T_177) begin
            if (4'hc == idxUpdate_4[3:0]) begin
              TBEAddr_12 <= 32'h0;
            end else begin
              TBEAddr_12 <= _GEN_2035;
            end
          end else begin
            TBEAddr_12 <= _GEN_2035;
          end
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEAddr_12 <= 32'h0;
          end else begin
            TBEAddr_12 <= _GEN_2549;
          end
        end else begin
          TBEAddr_12 <= _GEN_2549;
        end
      end else if (isAlloc_5) begin
        if (4'hc == idxAlloc[3:0]) begin
          TBEAddr_12 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_12 <= _GEN_2549;
        end
      end else if (_T_199) begin
        if (4'hc == idxUpdate_5[3:0]) begin
          TBEAddr_12 <= 32'h0;
        end else begin
          TBEAddr_12 <= _GEN_2549;
        end
      end else begin
        TBEAddr_12 <= _GEN_2549;
      end
    end else if (_T_243) begin
      if (4'hc == idxUpdate_7[3:0]) begin
        TBEAddr_12 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'hc == idxAlloc[3:0]) begin
          TBEAddr_12 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'hc == idxAlloc[3:0]) begin
            TBEAddr_12 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_12 <= _GEN_2549;
          end
        end else if (_T_199) begin
          if (4'hc == idxUpdate_5[3:0]) begin
            TBEAddr_12 <= 32'h0;
          end else begin
            TBEAddr_12 <= _GEN_2549;
          end
        end else begin
          TBEAddr_12 <= _GEN_2549;
        end
      end else if (_T_221) begin
        if (4'hc == idxUpdate_6[3:0]) begin
          TBEAddr_12 <= 32'h0;
        end else begin
          TBEAddr_12 <= _GEN_3063;
        end
      end else begin
        TBEAddr_12 <= _GEN_3063;
      end
    end else if (isAlloc_6) begin
      if (4'hc == idxAlloc[3:0]) begin
        TBEAddr_12 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_12 <= _GEN_3063;
      end
    end else if (_T_221) begin
      if (4'hc == idxUpdate_6[3:0]) begin
        TBEAddr_12 <= 32'h0;
      end else begin
        TBEAddr_12 <= _GEN_3063;
      end
    end else begin
      TBEAddr_12 <= _GEN_3063;
    end
    if (reset) begin
      TBEAddr_13 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'hd == idxAlloc[3:0]) begin
        TBEAddr_13 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'hd == idxAlloc[3:0]) begin
          TBEAddr_13 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEAddr_13 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEAddr_13 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEAddr_13 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEAddr_13 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEAddr_13 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEAddr_13 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEAddr_13 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEAddr_13 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEAddr_13 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEAddr_13 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEAddr_13 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'hd == idxUpdate_0[3:0]) begin
                    TBEAddr_13 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEAddr_13 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEAddr_13 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'hd == idxAlloc[3:0]) begin
                      TBEAddr_13 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'hd == idxUpdate_0[3:0]) begin
                      TBEAddr_13 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEAddr_13 <= 32'h0;
                  end else begin
                    TBEAddr_13 <= _GEN_494;
                  end
                end else begin
                  TBEAddr_13 <= _GEN_494;
                end
              end else if (isAlloc_1) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEAddr_13 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_13 <= _GEN_494;
                end
              end else if (_T_111) begin
                if (4'hd == idxUpdate_1[3:0]) begin
                  TBEAddr_13 <= 32'h0;
                end else begin
                  TBEAddr_13 <= _GEN_494;
                end
              end else begin
                TBEAddr_13 <= _GEN_494;
              end
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEAddr_13 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEAddr_13 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'hd == idxAlloc[3:0]) begin
                    TBEAddr_13 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_13 <= _GEN_494;
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUpdate_1[3:0]) begin
                    TBEAddr_13 <= 32'h0;
                  end else begin
                    TBEAddr_13 <= _GEN_494;
                  end
                end else begin
                  TBEAddr_13 <= _GEN_494;
                end
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEAddr_13 <= 32'h0;
                end else begin
                  TBEAddr_13 <= _GEN_1008;
                end
              end else begin
                TBEAddr_13 <= _GEN_1008;
              end
            end else if (isAlloc_2) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEAddr_13 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_13 <= _GEN_1008;
              end
            end else if (_T_133) begin
              if (4'hd == idxUpdate_2[3:0]) begin
                TBEAddr_13 <= 32'h0;
              end else begin
                TBEAddr_13 <= _GEN_1008;
              end
            end else begin
              TBEAddr_13 <= _GEN_1008;
            end
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEAddr_13 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEAddr_13 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'hd == idxAlloc[3:0]) begin
                  TBEAddr_13 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_13 <= _GEN_1008;
                end
              end else if (_T_133) begin
                if (4'hd == idxUpdate_2[3:0]) begin
                  TBEAddr_13 <= 32'h0;
                end else begin
                  TBEAddr_13 <= _GEN_1008;
                end
              end else begin
                TBEAddr_13 <= _GEN_1008;
              end
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEAddr_13 <= 32'h0;
              end else begin
                TBEAddr_13 <= _GEN_1522;
              end
            end else begin
              TBEAddr_13 <= _GEN_1522;
            end
          end else if (isAlloc_3) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEAddr_13 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_13 <= _GEN_1522;
            end
          end else if (_T_155) begin
            if (4'hd == idxUpdate_3[3:0]) begin
              TBEAddr_13 <= 32'h0;
            end else begin
              TBEAddr_13 <= _GEN_1522;
            end
          end else begin
            TBEAddr_13 <= _GEN_1522;
          end
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEAddr_13 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEAddr_13 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'hd == idxAlloc[3:0]) begin
                TBEAddr_13 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_13 <= _GEN_1522;
              end
            end else if (_T_155) begin
              if (4'hd == idxUpdate_3[3:0]) begin
                TBEAddr_13 <= 32'h0;
              end else begin
                TBEAddr_13 <= _GEN_1522;
              end
            end else begin
              TBEAddr_13 <= _GEN_1522;
            end
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEAddr_13 <= 32'h0;
            end else begin
              TBEAddr_13 <= _GEN_2036;
            end
          end else begin
            TBEAddr_13 <= _GEN_2036;
          end
        end else if (isAlloc_4) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEAddr_13 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_13 <= _GEN_2036;
          end
        end else if (_T_177) begin
          if (4'hd == idxUpdate_4[3:0]) begin
            TBEAddr_13 <= 32'h0;
          end else begin
            TBEAddr_13 <= _GEN_2036;
          end
        end else begin
          TBEAddr_13 <= _GEN_2036;
        end
      end else if (_T_221) begin
        if (4'hd == idxUpdate_6[3:0]) begin
          TBEAddr_13 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEAddr_13 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'hd == idxAlloc[3:0]) begin
              TBEAddr_13 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_13 <= _GEN_2036;
            end
          end else if (_T_177) begin
            if (4'hd == idxUpdate_4[3:0]) begin
              TBEAddr_13 <= 32'h0;
            end else begin
              TBEAddr_13 <= _GEN_2036;
            end
          end else begin
            TBEAddr_13 <= _GEN_2036;
          end
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEAddr_13 <= 32'h0;
          end else begin
            TBEAddr_13 <= _GEN_2550;
          end
        end else begin
          TBEAddr_13 <= _GEN_2550;
        end
      end else if (isAlloc_5) begin
        if (4'hd == idxAlloc[3:0]) begin
          TBEAddr_13 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_13 <= _GEN_2550;
        end
      end else if (_T_199) begin
        if (4'hd == idxUpdate_5[3:0]) begin
          TBEAddr_13 <= 32'h0;
        end else begin
          TBEAddr_13 <= _GEN_2550;
        end
      end else begin
        TBEAddr_13 <= _GEN_2550;
      end
    end else if (_T_243) begin
      if (4'hd == idxUpdate_7[3:0]) begin
        TBEAddr_13 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'hd == idxAlloc[3:0]) begin
          TBEAddr_13 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'hd == idxAlloc[3:0]) begin
            TBEAddr_13 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_13 <= _GEN_2550;
          end
        end else if (_T_199) begin
          if (4'hd == idxUpdate_5[3:0]) begin
            TBEAddr_13 <= 32'h0;
          end else begin
            TBEAddr_13 <= _GEN_2550;
          end
        end else begin
          TBEAddr_13 <= _GEN_2550;
        end
      end else if (_T_221) begin
        if (4'hd == idxUpdate_6[3:0]) begin
          TBEAddr_13 <= 32'h0;
        end else begin
          TBEAddr_13 <= _GEN_3064;
        end
      end else begin
        TBEAddr_13 <= _GEN_3064;
      end
    end else if (isAlloc_6) begin
      if (4'hd == idxAlloc[3:0]) begin
        TBEAddr_13 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_13 <= _GEN_3064;
      end
    end else if (_T_221) begin
      if (4'hd == idxUpdate_6[3:0]) begin
        TBEAddr_13 <= 32'h0;
      end else begin
        TBEAddr_13 <= _GEN_3064;
      end
    end else begin
      TBEAddr_13 <= _GEN_3064;
    end
    if (reset) begin
      TBEAddr_14 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'he == idxAlloc[3:0]) begin
        TBEAddr_14 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'he == idxAlloc[3:0]) begin
          TBEAddr_14 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEAddr_14 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEAddr_14 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEAddr_14 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEAddr_14 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEAddr_14 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEAddr_14 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEAddr_14 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEAddr_14 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEAddr_14 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEAddr_14 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEAddr_14 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'he == idxUpdate_0[3:0]) begin
                    TBEAddr_14 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEAddr_14 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEAddr_14 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'he == idxAlloc[3:0]) begin
                      TBEAddr_14 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'he == idxUpdate_0[3:0]) begin
                      TBEAddr_14 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEAddr_14 <= 32'h0;
                  end else begin
                    TBEAddr_14 <= _GEN_495;
                  end
                end else begin
                  TBEAddr_14 <= _GEN_495;
                end
              end else if (isAlloc_1) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEAddr_14 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_14 <= _GEN_495;
                end
              end else if (_T_111) begin
                if (4'he == idxUpdate_1[3:0]) begin
                  TBEAddr_14 <= 32'h0;
                end else begin
                  TBEAddr_14 <= _GEN_495;
                end
              end else begin
                TBEAddr_14 <= _GEN_495;
              end
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEAddr_14 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEAddr_14 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'he == idxAlloc[3:0]) begin
                    TBEAddr_14 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_14 <= _GEN_495;
                  end
                end else if (_T_111) begin
                  if (4'he == idxUpdate_1[3:0]) begin
                    TBEAddr_14 <= 32'h0;
                  end else begin
                    TBEAddr_14 <= _GEN_495;
                  end
                end else begin
                  TBEAddr_14 <= _GEN_495;
                end
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEAddr_14 <= 32'h0;
                end else begin
                  TBEAddr_14 <= _GEN_1009;
                end
              end else begin
                TBEAddr_14 <= _GEN_1009;
              end
            end else if (isAlloc_2) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEAddr_14 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_14 <= _GEN_1009;
              end
            end else if (_T_133) begin
              if (4'he == idxUpdate_2[3:0]) begin
                TBEAddr_14 <= 32'h0;
              end else begin
                TBEAddr_14 <= _GEN_1009;
              end
            end else begin
              TBEAddr_14 <= _GEN_1009;
            end
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEAddr_14 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEAddr_14 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'he == idxAlloc[3:0]) begin
                  TBEAddr_14 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_14 <= _GEN_1009;
                end
              end else if (_T_133) begin
                if (4'he == idxUpdate_2[3:0]) begin
                  TBEAddr_14 <= 32'h0;
                end else begin
                  TBEAddr_14 <= _GEN_1009;
                end
              end else begin
                TBEAddr_14 <= _GEN_1009;
              end
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEAddr_14 <= 32'h0;
              end else begin
                TBEAddr_14 <= _GEN_1523;
              end
            end else begin
              TBEAddr_14 <= _GEN_1523;
            end
          end else if (isAlloc_3) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEAddr_14 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_14 <= _GEN_1523;
            end
          end else if (_T_155) begin
            if (4'he == idxUpdate_3[3:0]) begin
              TBEAddr_14 <= 32'h0;
            end else begin
              TBEAddr_14 <= _GEN_1523;
            end
          end else begin
            TBEAddr_14 <= _GEN_1523;
          end
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEAddr_14 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEAddr_14 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'he == idxAlloc[3:0]) begin
                TBEAddr_14 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_14 <= _GEN_1523;
              end
            end else if (_T_155) begin
              if (4'he == idxUpdate_3[3:0]) begin
                TBEAddr_14 <= 32'h0;
              end else begin
                TBEAddr_14 <= _GEN_1523;
              end
            end else begin
              TBEAddr_14 <= _GEN_1523;
            end
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEAddr_14 <= 32'h0;
            end else begin
              TBEAddr_14 <= _GEN_2037;
            end
          end else begin
            TBEAddr_14 <= _GEN_2037;
          end
        end else if (isAlloc_4) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEAddr_14 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_14 <= _GEN_2037;
          end
        end else if (_T_177) begin
          if (4'he == idxUpdate_4[3:0]) begin
            TBEAddr_14 <= 32'h0;
          end else begin
            TBEAddr_14 <= _GEN_2037;
          end
        end else begin
          TBEAddr_14 <= _GEN_2037;
        end
      end else if (_T_221) begin
        if (4'he == idxUpdate_6[3:0]) begin
          TBEAddr_14 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEAddr_14 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'he == idxAlloc[3:0]) begin
              TBEAddr_14 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_14 <= _GEN_2037;
            end
          end else if (_T_177) begin
            if (4'he == idxUpdate_4[3:0]) begin
              TBEAddr_14 <= 32'h0;
            end else begin
              TBEAddr_14 <= _GEN_2037;
            end
          end else begin
            TBEAddr_14 <= _GEN_2037;
          end
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEAddr_14 <= 32'h0;
          end else begin
            TBEAddr_14 <= _GEN_2551;
          end
        end else begin
          TBEAddr_14 <= _GEN_2551;
        end
      end else if (isAlloc_5) begin
        if (4'he == idxAlloc[3:0]) begin
          TBEAddr_14 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_14 <= _GEN_2551;
        end
      end else if (_T_199) begin
        if (4'he == idxUpdate_5[3:0]) begin
          TBEAddr_14 <= 32'h0;
        end else begin
          TBEAddr_14 <= _GEN_2551;
        end
      end else begin
        TBEAddr_14 <= _GEN_2551;
      end
    end else if (_T_243) begin
      if (4'he == idxUpdate_7[3:0]) begin
        TBEAddr_14 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'he == idxAlloc[3:0]) begin
          TBEAddr_14 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'he == idxAlloc[3:0]) begin
            TBEAddr_14 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_14 <= _GEN_2551;
          end
        end else if (_T_199) begin
          if (4'he == idxUpdate_5[3:0]) begin
            TBEAddr_14 <= 32'h0;
          end else begin
            TBEAddr_14 <= _GEN_2551;
          end
        end else begin
          TBEAddr_14 <= _GEN_2551;
        end
      end else if (_T_221) begin
        if (4'he == idxUpdate_6[3:0]) begin
          TBEAddr_14 <= 32'h0;
        end else begin
          TBEAddr_14 <= _GEN_3065;
        end
      end else begin
        TBEAddr_14 <= _GEN_3065;
      end
    end else if (isAlloc_6) begin
      if (4'he == idxAlloc[3:0]) begin
        TBEAddr_14 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_14 <= _GEN_3065;
      end
    end else if (_T_221) begin
      if (4'he == idxUpdate_6[3:0]) begin
        TBEAddr_14 <= 32'h0;
      end else begin
        TBEAddr_14 <= _GEN_3065;
      end
    end else begin
      TBEAddr_14 <= _GEN_3065;
    end
    if (reset) begin
      TBEAddr_15 <= 32'h0;
    end else if (isAlloc_7) begin
      if (4'hf == idxAlloc[3:0]) begin
        TBEAddr_15 <= io_write_7_bits_addr[31:0];
      end else if (isAlloc_6) begin
        if (4'hf == idxAlloc[3:0]) begin
          TBEAddr_15 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEAddr_15 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEAddr_15 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEAddr_15 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEAddr_15 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEAddr_15 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEAddr_15 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEAddr_15 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEAddr_15 <= 32'h0;
                  end else if (isAlloc_0) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEAddr_15 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEAddr_15 <= 32'h0;
                    end
                  end
                end else if (isAlloc_0) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEAddr_15 <= io_write_0_bits_addr[31:0];
                  end
                end else if (_T_89) begin
                  if (4'hf == idxUpdate_0[3:0]) begin
                    TBEAddr_15 <= 32'h0;
                  end
                end
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEAddr_15 <= 32'h0;
                end else if (isAlloc_1) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEAddr_15 <= io_write_1_bits_addr[31:0];
                  end else if (isAlloc_0) begin
                    if (4'hf == idxAlloc[3:0]) begin
                      TBEAddr_15 <= io_write_0_bits_addr[31:0];
                    end
                  end else if (_T_89) begin
                    if (4'hf == idxUpdate_0[3:0]) begin
                      TBEAddr_15 <= 32'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEAddr_15 <= 32'h0;
                  end else begin
                    TBEAddr_15 <= _GEN_496;
                  end
                end else begin
                  TBEAddr_15 <= _GEN_496;
                end
              end else if (isAlloc_1) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEAddr_15 <= io_write_1_bits_addr[31:0];
                end else begin
                  TBEAddr_15 <= _GEN_496;
                end
              end else if (_T_111) begin
                if (4'hf == idxUpdate_1[3:0]) begin
                  TBEAddr_15 <= 32'h0;
                end else begin
                  TBEAddr_15 <= _GEN_496;
                end
              end else begin
                TBEAddr_15 <= _GEN_496;
              end
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEAddr_15 <= 32'h0;
              end else if (isAlloc_2) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEAddr_15 <= io_write_2_bits_addr[31:0];
                end else if (isAlloc_1) begin
                  if (4'hf == idxAlloc[3:0]) begin
                    TBEAddr_15 <= io_write_1_bits_addr[31:0];
                  end else begin
                    TBEAddr_15 <= _GEN_496;
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUpdate_1[3:0]) begin
                    TBEAddr_15 <= 32'h0;
                  end else begin
                    TBEAddr_15 <= _GEN_496;
                  end
                end else begin
                  TBEAddr_15 <= _GEN_496;
                end
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEAddr_15 <= 32'h0;
                end else begin
                  TBEAddr_15 <= _GEN_1010;
                end
              end else begin
                TBEAddr_15 <= _GEN_1010;
              end
            end else if (isAlloc_2) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEAddr_15 <= io_write_2_bits_addr[31:0];
              end else begin
                TBEAddr_15 <= _GEN_1010;
              end
            end else if (_T_133) begin
              if (4'hf == idxUpdate_2[3:0]) begin
                TBEAddr_15 <= 32'h0;
              end else begin
                TBEAddr_15 <= _GEN_1010;
              end
            end else begin
              TBEAddr_15 <= _GEN_1010;
            end
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEAddr_15 <= 32'h0;
            end else if (isAlloc_3) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEAddr_15 <= io_write_3_bits_addr[31:0];
              end else if (isAlloc_2) begin
                if (4'hf == idxAlloc[3:0]) begin
                  TBEAddr_15 <= io_write_2_bits_addr[31:0];
                end else begin
                  TBEAddr_15 <= _GEN_1010;
                end
              end else if (_T_133) begin
                if (4'hf == idxUpdate_2[3:0]) begin
                  TBEAddr_15 <= 32'h0;
                end else begin
                  TBEAddr_15 <= _GEN_1010;
                end
              end else begin
                TBEAddr_15 <= _GEN_1010;
              end
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEAddr_15 <= 32'h0;
              end else begin
                TBEAddr_15 <= _GEN_1524;
              end
            end else begin
              TBEAddr_15 <= _GEN_1524;
            end
          end else if (isAlloc_3) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEAddr_15 <= io_write_3_bits_addr[31:0];
            end else begin
              TBEAddr_15 <= _GEN_1524;
            end
          end else if (_T_155) begin
            if (4'hf == idxUpdate_3[3:0]) begin
              TBEAddr_15 <= 32'h0;
            end else begin
              TBEAddr_15 <= _GEN_1524;
            end
          end else begin
            TBEAddr_15 <= _GEN_1524;
          end
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEAddr_15 <= 32'h0;
          end else if (isAlloc_4) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEAddr_15 <= io_write_4_bits_addr[31:0];
            end else if (isAlloc_3) begin
              if (4'hf == idxAlloc[3:0]) begin
                TBEAddr_15 <= io_write_3_bits_addr[31:0];
              end else begin
                TBEAddr_15 <= _GEN_1524;
              end
            end else if (_T_155) begin
              if (4'hf == idxUpdate_3[3:0]) begin
                TBEAddr_15 <= 32'h0;
              end else begin
                TBEAddr_15 <= _GEN_1524;
              end
            end else begin
              TBEAddr_15 <= _GEN_1524;
            end
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEAddr_15 <= 32'h0;
            end else begin
              TBEAddr_15 <= _GEN_2038;
            end
          end else begin
            TBEAddr_15 <= _GEN_2038;
          end
        end else if (isAlloc_4) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEAddr_15 <= io_write_4_bits_addr[31:0];
          end else begin
            TBEAddr_15 <= _GEN_2038;
          end
        end else if (_T_177) begin
          if (4'hf == idxUpdate_4[3:0]) begin
            TBEAddr_15 <= 32'h0;
          end else begin
            TBEAddr_15 <= _GEN_2038;
          end
        end else begin
          TBEAddr_15 <= _GEN_2038;
        end
      end else if (_T_221) begin
        if (4'hf == idxUpdate_6[3:0]) begin
          TBEAddr_15 <= 32'h0;
        end else if (isAlloc_5) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEAddr_15 <= io_write_5_bits_addr[31:0];
          end else if (isAlloc_4) begin
            if (4'hf == idxAlloc[3:0]) begin
              TBEAddr_15 <= io_write_4_bits_addr[31:0];
            end else begin
              TBEAddr_15 <= _GEN_2038;
            end
          end else if (_T_177) begin
            if (4'hf == idxUpdate_4[3:0]) begin
              TBEAddr_15 <= 32'h0;
            end else begin
              TBEAddr_15 <= _GEN_2038;
            end
          end else begin
            TBEAddr_15 <= _GEN_2038;
          end
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEAddr_15 <= 32'h0;
          end else begin
            TBEAddr_15 <= _GEN_2552;
          end
        end else begin
          TBEAddr_15 <= _GEN_2552;
        end
      end else if (isAlloc_5) begin
        if (4'hf == idxAlloc[3:0]) begin
          TBEAddr_15 <= io_write_5_bits_addr[31:0];
        end else begin
          TBEAddr_15 <= _GEN_2552;
        end
      end else if (_T_199) begin
        if (4'hf == idxUpdate_5[3:0]) begin
          TBEAddr_15 <= 32'h0;
        end else begin
          TBEAddr_15 <= _GEN_2552;
        end
      end else begin
        TBEAddr_15 <= _GEN_2552;
      end
    end else if (_T_243) begin
      if (4'hf == idxUpdate_7[3:0]) begin
        TBEAddr_15 <= 32'h0;
      end else if (isAlloc_6) begin
        if (4'hf == idxAlloc[3:0]) begin
          TBEAddr_15 <= io_write_6_bits_addr[31:0];
        end else if (isAlloc_5) begin
          if (4'hf == idxAlloc[3:0]) begin
            TBEAddr_15 <= io_write_5_bits_addr[31:0];
          end else begin
            TBEAddr_15 <= _GEN_2552;
          end
        end else if (_T_199) begin
          if (4'hf == idxUpdate_5[3:0]) begin
            TBEAddr_15 <= 32'h0;
          end else begin
            TBEAddr_15 <= _GEN_2552;
          end
        end else begin
          TBEAddr_15 <= _GEN_2552;
        end
      end else if (_T_221) begin
        if (4'hf == idxUpdate_6[3:0]) begin
          TBEAddr_15 <= 32'h0;
        end else begin
          TBEAddr_15 <= _GEN_3066;
        end
      end else begin
        TBEAddr_15 <= _GEN_3066;
      end
    end else if (isAlloc_6) begin
      if (4'hf == idxAlloc[3:0]) begin
        TBEAddr_15 <= io_write_6_bits_addr[31:0];
      end else begin
        TBEAddr_15 <= _GEN_3066;
      end
    end else if (_T_221) begin
      if (4'hf == idxUpdate_6[3:0]) begin
        TBEAddr_15 <= 32'h0;
      end else begin
        TBEAddr_15 <= _GEN_3066;
      end
    end else begin
      TBEAddr_15 <= _GEN_3066;
    end
    if (reset) begin
      counter <= 6'h0;
    end else if (isAlloc_7) begin
      counter <= _T_88;
    end else if (_T_243) begin
      counter <= _T_96;
    end else if (isAlloc_6) begin
      counter <= _T_88;
    end else if (_T_221) begin
      counter <= _T_96;
    end else if (isAlloc_5) begin
      counter <= _T_88;
    end else if (_T_199) begin
      counter <= _T_96;
    end else if (isAlloc_4) begin
      counter <= _T_88;
    end else if (_T_177) begin
      counter <= _T_96;
    end else if (isAlloc_3) begin
      counter <= _T_88;
    end else if (_T_155) begin
      counter <= _T_96;
    end else if (isAlloc_2) begin
      counter <= _T_88;
    end else if (_T_133) begin
      counter <= _T_96;
    end else if (isAlloc_1) begin
      counter <= _T_88;
    end else if (_T_111) begin
      counter <= _T_96;
    end else if (isAlloc_0) begin
      counter <= _T_88;
    end else if (_T_89) begin
      counter <= _T_96;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_4293 & _T_102) begin
          $fwrite(32'h80000002,"TBE Field Check %d\n",_GEN_223); // @[TBE.scala 122:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_4298 & _T_102) begin
          $fwrite(32'h80000002,"TBE Field Check %d\n",_GEN_737); // @[TBE.scala 122:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_4303 & _T_102) begin
          $fwrite(32'h80000002,"TBE Field Check %d\n",_GEN_1251); // @[TBE.scala 122:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_4308 & _T_102) begin
          $fwrite(32'h80000002,"TBE Field Check %d\n",_GEN_1765); // @[TBE.scala 122:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_4313 & _T_102) begin
          $fwrite(32'h80000002,"TBE Field Check %d\n",_GEN_2279); // @[TBE.scala 122:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_4318 & _T_102) begin
          $fwrite(32'h80000002,"TBE Field Check %d\n",_GEN_2793); // @[TBE.scala 122:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_4323 & _T_102) begin
          $fwrite(32'h80000002,"TBE Field Check %d\n",_GEN_3307); // @[TBE.scala 122:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_4328 & _T_102) begin
          $fwrite(32'h80000002,"TBE Field Check %d\n",_GEN_3821); // @[TBE.scala 122:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module lockVector(
  input         clock,
  input         reset,
  input         io_lock_in_valid,
  input  [31:0] io_lock_in_bits_addr,
  output        io_probe_out_valid,
  output        io_probe_out_bits,
  input         io_probe_in_valid,
  input  [31:0] io_probe_in_bits_addr,
  input         io_unLock_0_in_valid,
  input  [31:0] io_unLock_0_in_bits_addr,
  input         io_unLock_1_in_valid,
  input  [31:0] io_unLock_1_in_bits_addr,
  input         io_unLock_2_in_valid,
  input  [31:0] io_unLock_2_in_bits_addr,
  input         io_unLock_3_in_valid,
  input  [31:0] io_unLock_3_in_bits_addr,
  input         io_unLock_4_in_valid,
  input  [31:0] io_unLock_4_in_bits_addr,
  input         io_unLock_5_in_valid,
  input  [31:0] io_unLock_5_in_bits_addr,
  input         io_unLock_6_in_valid,
  input  [31:0] io_unLock_6_in_bits_addr,
  input         io_unLock_7_in_valid,
  input  [31:0] io_unLock_7_in_bits_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] finder_0_io_key; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_0; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_1; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_2; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_3; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_4; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_5; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_6; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_7; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_8; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_9; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_10; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_11; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_12; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_13; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_14; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_15; // @[elements.scala 158:28]
  wire  finder_0_io_valid_0; // @[elements.scala 158:28]
  wire  finder_0_io_valid_1; // @[elements.scala 158:28]
  wire  finder_0_io_valid_2; // @[elements.scala 158:28]
  wire  finder_0_io_valid_3; // @[elements.scala 158:28]
  wire  finder_0_io_valid_4; // @[elements.scala 158:28]
  wire  finder_0_io_valid_5; // @[elements.scala 158:28]
  wire  finder_0_io_valid_6; // @[elements.scala 158:28]
  wire  finder_0_io_valid_7; // @[elements.scala 158:28]
  wire  finder_0_io_valid_8; // @[elements.scala 158:28]
  wire  finder_0_io_valid_9; // @[elements.scala 158:28]
  wire  finder_0_io_valid_10; // @[elements.scala 158:28]
  wire  finder_0_io_valid_11; // @[elements.scala 158:28]
  wire  finder_0_io_valid_12; // @[elements.scala 158:28]
  wire  finder_0_io_valid_13; // @[elements.scala 158:28]
  wire  finder_0_io_valid_14; // @[elements.scala 158:28]
  wire  finder_0_io_valid_15; // @[elements.scala 158:28]
  wire  finder_0_io_value_valid; // @[elements.scala 158:28]
  wire [3:0] finder_0_io_value_bits; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_key; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_0; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_1; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_2; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_3; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_4; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_5; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_6; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_7; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_8; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_9; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_10; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_11; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_12; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_13; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_14; // @[elements.scala 158:28]
  wire [31:0] finder_1_io_data_15; // @[elements.scala 158:28]
  wire  finder_1_io_valid_0; // @[elements.scala 158:28]
  wire  finder_1_io_valid_1; // @[elements.scala 158:28]
  wire  finder_1_io_valid_2; // @[elements.scala 158:28]
  wire  finder_1_io_valid_3; // @[elements.scala 158:28]
  wire  finder_1_io_valid_4; // @[elements.scala 158:28]
  wire  finder_1_io_valid_5; // @[elements.scala 158:28]
  wire  finder_1_io_valid_6; // @[elements.scala 158:28]
  wire  finder_1_io_valid_7; // @[elements.scala 158:28]
  wire  finder_1_io_valid_8; // @[elements.scala 158:28]
  wire  finder_1_io_valid_9; // @[elements.scala 158:28]
  wire  finder_1_io_valid_10; // @[elements.scala 158:28]
  wire  finder_1_io_valid_11; // @[elements.scala 158:28]
  wire  finder_1_io_valid_12; // @[elements.scala 158:28]
  wire  finder_1_io_valid_13; // @[elements.scala 158:28]
  wire  finder_1_io_valid_14; // @[elements.scala 158:28]
  wire  finder_1_io_valid_15; // @[elements.scala 158:28]
  wire  finder_1_io_value_valid; // @[elements.scala 158:28]
  wire [3:0] finder_1_io_value_bits; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_key; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_0; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_1; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_2; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_3; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_4; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_5; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_6; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_7; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_8; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_9; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_10; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_11; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_12; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_13; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_14; // @[elements.scala 158:28]
  wire [31:0] finder_2_io_data_15; // @[elements.scala 158:28]
  wire  finder_2_io_valid_0; // @[elements.scala 158:28]
  wire  finder_2_io_valid_1; // @[elements.scala 158:28]
  wire  finder_2_io_valid_2; // @[elements.scala 158:28]
  wire  finder_2_io_valid_3; // @[elements.scala 158:28]
  wire  finder_2_io_valid_4; // @[elements.scala 158:28]
  wire  finder_2_io_valid_5; // @[elements.scala 158:28]
  wire  finder_2_io_valid_6; // @[elements.scala 158:28]
  wire  finder_2_io_valid_7; // @[elements.scala 158:28]
  wire  finder_2_io_valid_8; // @[elements.scala 158:28]
  wire  finder_2_io_valid_9; // @[elements.scala 158:28]
  wire  finder_2_io_valid_10; // @[elements.scala 158:28]
  wire  finder_2_io_valid_11; // @[elements.scala 158:28]
  wire  finder_2_io_valid_12; // @[elements.scala 158:28]
  wire  finder_2_io_valid_13; // @[elements.scala 158:28]
  wire  finder_2_io_valid_14; // @[elements.scala 158:28]
  wire  finder_2_io_valid_15; // @[elements.scala 158:28]
  wire  finder_2_io_value_valid; // @[elements.scala 158:28]
  wire [3:0] finder_2_io_value_bits; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_key; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_0; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_1; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_2; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_3; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_4; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_5; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_6; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_7; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_8; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_9; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_10; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_11; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_12; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_13; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_14; // @[elements.scala 158:28]
  wire [31:0] finder_3_io_data_15; // @[elements.scala 158:28]
  wire  finder_3_io_valid_0; // @[elements.scala 158:28]
  wire  finder_3_io_valid_1; // @[elements.scala 158:28]
  wire  finder_3_io_valid_2; // @[elements.scala 158:28]
  wire  finder_3_io_valid_3; // @[elements.scala 158:28]
  wire  finder_3_io_valid_4; // @[elements.scala 158:28]
  wire  finder_3_io_valid_5; // @[elements.scala 158:28]
  wire  finder_3_io_valid_6; // @[elements.scala 158:28]
  wire  finder_3_io_valid_7; // @[elements.scala 158:28]
  wire  finder_3_io_valid_8; // @[elements.scala 158:28]
  wire  finder_3_io_valid_9; // @[elements.scala 158:28]
  wire  finder_3_io_valid_10; // @[elements.scala 158:28]
  wire  finder_3_io_valid_11; // @[elements.scala 158:28]
  wire  finder_3_io_valid_12; // @[elements.scala 158:28]
  wire  finder_3_io_valid_13; // @[elements.scala 158:28]
  wire  finder_3_io_valid_14; // @[elements.scala 158:28]
  wire  finder_3_io_valid_15; // @[elements.scala 158:28]
  wire  finder_3_io_value_valid; // @[elements.scala 158:28]
  wire [3:0] finder_3_io_value_bits; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_key; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_0; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_1; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_2; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_3; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_4; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_5; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_6; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_7; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_8; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_9; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_10; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_11; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_12; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_13; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_14; // @[elements.scala 158:28]
  wire [31:0] finder_4_io_data_15; // @[elements.scala 158:28]
  wire  finder_4_io_valid_0; // @[elements.scala 158:28]
  wire  finder_4_io_valid_1; // @[elements.scala 158:28]
  wire  finder_4_io_valid_2; // @[elements.scala 158:28]
  wire  finder_4_io_valid_3; // @[elements.scala 158:28]
  wire  finder_4_io_valid_4; // @[elements.scala 158:28]
  wire  finder_4_io_valid_5; // @[elements.scala 158:28]
  wire  finder_4_io_valid_6; // @[elements.scala 158:28]
  wire  finder_4_io_valid_7; // @[elements.scala 158:28]
  wire  finder_4_io_valid_8; // @[elements.scala 158:28]
  wire  finder_4_io_valid_9; // @[elements.scala 158:28]
  wire  finder_4_io_valid_10; // @[elements.scala 158:28]
  wire  finder_4_io_valid_11; // @[elements.scala 158:28]
  wire  finder_4_io_valid_12; // @[elements.scala 158:28]
  wire  finder_4_io_valid_13; // @[elements.scala 158:28]
  wire  finder_4_io_valid_14; // @[elements.scala 158:28]
  wire  finder_4_io_valid_15; // @[elements.scala 158:28]
  wire  finder_4_io_value_valid; // @[elements.scala 158:28]
  wire [3:0] finder_4_io_value_bits; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_key; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_0; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_1; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_2; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_3; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_4; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_5; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_6; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_7; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_8; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_9; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_10; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_11; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_12; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_13; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_14; // @[elements.scala 158:28]
  wire [31:0] finder_5_io_data_15; // @[elements.scala 158:28]
  wire  finder_5_io_valid_0; // @[elements.scala 158:28]
  wire  finder_5_io_valid_1; // @[elements.scala 158:28]
  wire  finder_5_io_valid_2; // @[elements.scala 158:28]
  wire  finder_5_io_valid_3; // @[elements.scala 158:28]
  wire  finder_5_io_valid_4; // @[elements.scala 158:28]
  wire  finder_5_io_valid_5; // @[elements.scala 158:28]
  wire  finder_5_io_valid_6; // @[elements.scala 158:28]
  wire  finder_5_io_valid_7; // @[elements.scala 158:28]
  wire  finder_5_io_valid_8; // @[elements.scala 158:28]
  wire  finder_5_io_valid_9; // @[elements.scala 158:28]
  wire  finder_5_io_valid_10; // @[elements.scala 158:28]
  wire  finder_5_io_valid_11; // @[elements.scala 158:28]
  wire  finder_5_io_valid_12; // @[elements.scala 158:28]
  wire  finder_5_io_valid_13; // @[elements.scala 158:28]
  wire  finder_5_io_valid_14; // @[elements.scala 158:28]
  wire  finder_5_io_valid_15; // @[elements.scala 158:28]
  wire  finder_5_io_value_valid; // @[elements.scala 158:28]
  wire [3:0] finder_5_io_value_bits; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_key; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_0; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_1; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_2; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_3; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_4; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_5; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_6; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_7; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_8; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_9; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_10; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_11; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_12; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_13; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_14; // @[elements.scala 158:28]
  wire [31:0] finder_6_io_data_15; // @[elements.scala 158:28]
  wire  finder_6_io_valid_0; // @[elements.scala 158:28]
  wire  finder_6_io_valid_1; // @[elements.scala 158:28]
  wire  finder_6_io_valid_2; // @[elements.scala 158:28]
  wire  finder_6_io_valid_3; // @[elements.scala 158:28]
  wire  finder_6_io_valid_4; // @[elements.scala 158:28]
  wire  finder_6_io_valid_5; // @[elements.scala 158:28]
  wire  finder_6_io_valid_6; // @[elements.scala 158:28]
  wire  finder_6_io_valid_7; // @[elements.scala 158:28]
  wire  finder_6_io_valid_8; // @[elements.scala 158:28]
  wire  finder_6_io_valid_9; // @[elements.scala 158:28]
  wire  finder_6_io_valid_10; // @[elements.scala 158:28]
  wire  finder_6_io_valid_11; // @[elements.scala 158:28]
  wire  finder_6_io_valid_12; // @[elements.scala 158:28]
  wire  finder_6_io_valid_13; // @[elements.scala 158:28]
  wire  finder_6_io_valid_14; // @[elements.scala 158:28]
  wire  finder_6_io_valid_15; // @[elements.scala 158:28]
  wire  finder_6_io_value_valid; // @[elements.scala 158:28]
  wire [3:0] finder_6_io_value_bits; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_key; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_0; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_1; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_2; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_3; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_4; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_5; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_6; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_7; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_8; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_9; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_10; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_11; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_12; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_13; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_14; // @[elements.scala 158:28]
  wire [31:0] finder_7_io_data_15; // @[elements.scala 158:28]
  wire  finder_7_io_valid_0; // @[elements.scala 158:28]
  wire  finder_7_io_valid_1; // @[elements.scala 158:28]
  wire  finder_7_io_valid_2; // @[elements.scala 158:28]
  wire  finder_7_io_valid_3; // @[elements.scala 158:28]
  wire  finder_7_io_valid_4; // @[elements.scala 158:28]
  wire  finder_7_io_valid_5; // @[elements.scala 158:28]
  wire  finder_7_io_valid_6; // @[elements.scala 158:28]
  wire  finder_7_io_valid_7; // @[elements.scala 158:28]
  wire  finder_7_io_valid_8; // @[elements.scala 158:28]
  wire  finder_7_io_valid_9; // @[elements.scala 158:28]
  wire  finder_7_io_valid_10; // @[elements.scala 158:28]
  wire  finder_7_io_valid_11; // @[elements.scala 158:28]
  wire  finder_7_io_valid_12; // @[elements.scala 158:28]
  wire  finder_7_io_valid_13; // @[elements.scala 158:28]
  wire  finder_7_io_valid_14; // @[elements.scala 158:28]
  wire  finder_7_io_valid_15; // @[elements.scala 158:28]
  wire  finder_7_io_value_valid; // @[elements.scala 158:28]
  wire [3:0] finder_7_io_value_bits; // @[elements.scala 158:28]
  reg [31:0] addrVec_0; // @[elements.scala 148:26]
  reg [31:0] addrVec_1; // @[elements.scala 148:26]
  reg [31:0] addrVec_2; // @[elements.scala 148:26]
  reg [31:0] addrVec_3; // @[elements.scala 148:26]
  reg [31:0] addrVec_4; // @[elements.scala 148:26]
  reg [31:0] addrVec_5; // @[elements.scala 148:26]
  reg [31:0] addrVec_6; // @[elements.scala 148:26]
  reg [31:0] addrVec_7; // @[elements.scala 148:26]
  reg [31:0] addrVec_8; // @[elements.scala 148:26]
  reg [31:0] addrVec_9; // @[elements.scala 148:26]
  reg [31:0] addrVec_10; // @[elements.scala 148:26]
  reg [31:0] addrVec_11; // @[elements.scala 148:26]
  reg [31:0] addrVec_12; // @[elements.scala 148:26]
  reg [31:0] addrVec_13; // @[elements.scala 148:26]
  reg [31:0] addrVec_14; // @[elements.scala 148:26]
  reg [31:0] addrVec_15; // @[elements.scala 148:26]
  reg  valid_0; // @[elements.scala 149:26]
  reg  valid_1; // @[elements.scala 149:26]
  reg  valid_2; // @[elements.scala 149:26]
  reg  valid_3; // @[elements.scala 149:26]
  reg  valid_4; // @[elements.scala 149:26]
  reg  valid_5; // @[elements.scala 149:26]
  reg  valid_6; // @[elements.scala 149:26]
  reg  valid_7; // @[elements.scala 149:26]
  reg  valid_8; // @[elements.scala 149:26]
  reg  valid_9; // @[elements.scala 149:26]
  reg  valid_10; // @[elements.scala 149:26]
  reg  valid_11; // @[elements.scala 149:26]
  reg  valid_12; // @[elements.scala 149:26]
  reg  valid_13; // @[elements.scala 149:26]
  reg  valid_14; // @[elements.scala 149:26]
  reg  valid_15; // @[elements.scala 149:26]
  wire  _T_39 = addrVec_15 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_37 = addrVec_14 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_35 = addrVec_13 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_33 = addrVec_12 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_31 = addrVec_11 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_29 = addrVec_10 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_27 = addrVec_9 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_25 = addrVec_8 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_23 = addrVec_7 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_21 = addrVec_6 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_19 = addrVec_5 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_17 = addrVec_4 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_15 = addrVec_3 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_13 = addrVec_2 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_11 = addrVec_1 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire  _T_9 = addrVec_0 == io_probe_in_bits_addr; // @[elements.scala 175:53]
  wire [7:0] _T_46 = {_T_23,_T_21,_T_19,_T_17,_T_15,_T_13,_T_11,_T_9}; // @[Cat.scala 29:58]
  wire [15:0] bitmapProbe = {_T_39,_T_37,_T_35,_T_33,_T_31,_T_29,_T_27,_T_25,_T_46}; // @[Cat.scala 29:58]
  wire [7:0] _T_149 = {valid_7,valid_6,valid_5,valid_4,valid_3,valid_2,valid_1,valid_0}; // @[elements.scala 201:45]
  wire [15:0] _T_157 = {valid_15,valid_14,valid_13,valid_12,valid_11,valid_10,valid_9,valid_8,_T_149}; // @[elements.scala 201:45]
  wire [15:0] _T_158 = bitmapProbe & _T_157; // @[elements.scala 201:31]
  wire  isLocked = _T_158 != 16'h0; // @[elements.scala 201:49]
  wire  _T_4 = ~isLocked; // @[elements.scala 171:28]
  wire  write = _T_4 & io_lock_in_valid; // @[elements.scala 171:38]
  wire  _T_111 = io_unLock_0_in_valid & finder_0_io_value_valid; // @[elements.scala 189:23]
  wire [15:0] idxUnlock_0 = {{12'd0}, finder_0_io_value_bits}; // @[elements.scala 155:26 elements.scala 185:22]
  wire  _GEN_0 = 4'h0 == idxUnlock_0[3:0] ? 1'h0 : valid_0; // @[elements.scala 190:33]
  wire  _GEN_1 = 4'h1 == idxUnlock_0[3:0] ? 1'h0 : valid_1; // @[elements.scala 190:33]
  wire  _GEN_2 = 4'h2 == idxUnlock_0[3:0] ? 1'h0 : valid_2; // @[elements.scala 190:33]
  wire  _GEN_3 = 4'h3 == idxUnlock_0[3:0] ? 1'h0 : valid_3; // @[elements.scala 190:33]
  wire  _GEN_4 = 4'h4 == idxUnlock_0[3:0] ? 1'h0 : valid_4; // @[elements.scala 190:33]
  wire  _GEN_5 = 4'h5 == idxUnlock_0[3:0] ? 1'h0 : valid_5; // @[elements.scala 190:33]
  wire  _GEN_6 = 4'h6 == idxUnlock_0[3:0] ? 1'h0 : valid_6; // @[elements.scala 190:33]
  wire  _GEN_7 = 4'h7 == idxUnlock_0[3:0] ? 1'h0 : valid_7; // @[elements.scala 190:33]
  wire  _GEN_8 = 4'h8 == idxUnlock_0[3:0] ? 1'h0 : valid_8; // @[elements.scala 190:33]
  wire  _GEN_9 = 4'h9 == idxUnlock_0[3:0] ? 1'h0 : valid_9; // @[elements.scala 190:33]
  wire  _GEN_10 = 4'ha == idxUnlock_0[3:0] ? 1'h0 : valid_10; // @[elements.scala 190:33]
  wire  _GEN_11 = 4'hb == idxUnlock_0[3:0] ? 1'h0 : valid_11; // @[elements.scala 190:33]
  wire  _GEN_12 = 4'hc == idxUnlock_0[3:0] ? 1'h0 : valid_12; // @[elements.scala 190:33]
  wire  _GEN_13 = 4'hd == idxUnlock_0[3:0] ? 1'h0 : valid_13; // @[elements.scala 190:33]
  wire  _GEN_14 = 4'he == idxUnlock_0[3:0] ? 1'h0 : valid_14; // @[elements.scala 190:33]
  wire  _GEN_15 = 4'hf == idxUnlock_0[3:0] ? 1'h0 : valid_15; // @[elements.scala 190:33]
  wire  _GEN_16 = _T_111 ? _GEN_0 : valid_0; // @[elements.scala 189:52]
  wire  _GEN_17 = _T_111 ? _GEN_1 : valid_1; // @[elements.scala 189:52]
  wire  _GEN_18 = _T_111 ? _GEN_2 : valid_2; // @[elements.scala 189:52]
  wire  _GEN_19 = _T_111 ? _GEN_3 : valid_3; // @[elements.scala 189:52]
  wire  _GEN_20 = _T_111 ? _GEN_4 : valid_4; // @[elements.scala 189:52]
  wire  _GEN_21 = _T_111 ? _GEN_5 : valid_5; // @[elements.scala 189:52]
  wire  _GEN_22 = _T_111 ? _GEN_6 : valid_6; // @[elements.scala 189:52]
  wire  _GEN_23 = _T_111 ? _GEN_7 : valid_7; // @[elements.scala 189:52]
  wire  _GEN_24 = _T_111 ? _GEN_8 : valid_8; // @[elements.scala 189:52]
  wire  _GEN_25 = _T_111 ? _GEN_9 : valid_9; // @[elements.scala 189:52]
  wire  _GEN_26 = _T_111 ? _GEN_10 : valid_10; // @[elements.scala 189:52]
  wire  _GEN_27 = _T_111 ? _GEN_11 : valid_11; // @[elements.scala 189:52]
  wire  _GEN_28 = _T_111 ? _GEN_12 : valid_12; // @[elements.scala 189:52]
  wire  _GEN_29 = _T_111 ? _GEN_13 : valid_13; // @[elements.scala 189:52]
  wire  _GEN_30 = _T_111 ? _GEN_14 : valid_14; // @[elements.scala 189:52]
  wire  _GEN_31 = _T_111 ? _GEN_15 : valid_15; // @[elements.scala 189:52]
  wire  _T_113 = io_unLock_1_in_valid & finder_1_io_value_valid; // @[elements.scala 189:23]
  wire [15:0] idxUnlock_1 = {{12'd0}, finder_1_io_value_bits}; // @[elements.scala 155:26 elements.scala 185:22]
  wire  _GEN_32 = 4'h0 == idxUnlock_1[3:0] ? 1'h0 : _GEN_16; // @[elements.scala 190:33]
  wire  _GEN_33 = 4'h1 == idxUnlock_1[3:0] ? 1'h0 : _GEN_17; // @[elements.scala 190:33]
  wire  _GEN_34 = 4'h2 == idxUnlock_1[3:0] ? 1'h0 : _GEN_18; // @[elements.scala 190:33]
  wire  _GEN_35 = 4'h3 == idxUnlock_1[3:0] ? 1'h0 : _GEN_19; // @[elements.scala 190:33]
  wire  _GEN_36 = 4'h4 == idxUnlock_1[3:0] ? 1'h0 : _GEN_20; // @[elements.scala 190:33]
  wire  _GEN_37 = 4'h5 == idxUnlock_1[3:0] ? 1'h0 : _GEN_21; // @[elements.scala 190:33]
  wire  _GEN_38 = 4'h6 == idxUnlock_1[3:0] ? 1'h0 : _GEN_22; // @[elements.scala 190:33]
  wire  _GEN_39 = 4'h7 == idxUnlock_1[3:0] ? 1'h0 : _GEN_23; // @[elements.scala 190:33]
  wire  _GEN_40 = 4'h8 == idxUnlock_1[3:0] ? 1'h0 : _GEN_24; // @[elements.scala 190:33]
  wire  _GEN_41 = 4'h9 == idxUnlock_1[3:0] ? 1'h0 : _GEN_25; // @[elements.scala 190:33]
  wire  _GEN_42 = 4'ha == idxUnlock_1[3:0] ? 1'h0 : _GEN_26; // @[elements.scala 190:33]
  wire  _GEN_43 = 4'hb == idxUnlock_1[3:0] ? 1'h0 : _GEN_27; // @[elements.scala 190:33]
  wire  _GEN_44 = 4'hc == idxUnlock_1[3:0] ? 1'h0 : _GEN_28; // @[elements.scala 190:33]
  wire  _GEN_45 = 4'hd == idxUnlock_1[3:0] ? 1'h0 : _GEN_29; // @[elements.scala 190:33]
  wire  _GEN_46 = 4'he == idxUnlock_1[3:0] ? 1'h0 : _GEN_30; // @[elements.scala 190:33]
  wire  _GEN_47 = 4'hf == idxUnlock_1[3:0] ? 1'h0 : _GEN_31; // @[elements.scala 190:33]
  wire  _GEN_48 = _T_113 ? _GEN_32 : _GEN_16; // @[elements.scala 189:52]
  wire  _GEN_49 = _T_113 ? _GEN_33 : _GEN_17; // @[elements.scala 189:52]
  wire  _GEN_50 = _T_113 ? _GEN_34 : _GEN_18; // @[elements.scala 189:52]
  wire  _GEN_51 = _T_113 ? _GEN_35 : _GEN_19; // @[elements.scala 189:52]
  wire  _GEN_52 = _T_113 ? _GEN_36 : _GEN_20; // @[elements.scala 189:52]
  wire  _GEN_53 = _T_113 ? _GEN_37 : _GEN_21; // @[elements.scala 189:52]
  wire  _GEN_54 = _T_113 ? _GEN_38 : _GEN_22; // @[elements.scala 189:52]
  wire  _GEN_55 = _T_113 ? _GEN_39 : _GEN_23; // @[elements.scala 189:52]
  wire  _GEN_56 = _T_113 ? _GEN_40 : _GEN_24; // @[elements.scala 189:52]
  wire  _GEN_57 = _T_113 ? _GEN_41 : _GEN_25; // @[elements.scala 189:52]
  wire  _GEN_58 = _T_113 ? _GEN_42 : _GEN_26; // @[elements.scala 189:52]
  wire  _GEN_59 = _T_113 ? _GEN_43 : _GEN_27; // @[elements.scala 189:52]
  wire  _GEN_60 = _T_113 ? _GEN_44 : _GEN_28; // @[elements.scala 189:52]
  wire  _GEN_61 = _T_113 ? _GEN_45 : _GEN_29; // @[elements.scala 189:52]
  wire  _GEN_62 = _T_113 ? _GEN_46 : _GEN_30; // @[elements.scala 189:52]
  wire  _GEN_63 = _T_113 ? _GEN_47 : _GEN_31; // @[elements.scala 189:52]
  wire  _T_115 = io_unLock_2_in_valid & finder_2_io_value_valid; // @[elements.scala 189:23]
  wire [15:0] idxUnlock_2 = {{12'd0}, finder_2_io_value_bits}; // @[elements.scala 155:26 elements.scala 185:22]
  wire  _GEN_64 = 4'h0 == idxUnlock_2[3:0] ? 1'h0 : _GEN_48; // @[elements.scala 190:33]
  wire  _GEN_65 = 4'h1 == idxUnlock_2[3:0] ? 1'h0 : _GEN_49; // @[elements.scala 190:33]
  wire  _GEN_66 = 4'h2 == idxUnlock_2[3:0] ? 1'h0 : _GEN_50; // @[elements.scala 190:33]
  wire  _GEN_67 = 4'h3 == idxUnlock_2[3:0] ? 1'h0 : _GEN_51; // @[elements.scala 190:33]
  wire  _GEN_68 = 4'h4 == idxUnlock_2[3:0] ? 1'h0 : _GEN_52; // @[elements.scala 190:33]
  wire  _GEN_69 = 4'h5 == idxUnlock_2[3:0] ? 1'h0 : _GEN_53; // @[elements.scala 190:33]
  wire  _GEN_70 = 4'h6 == idxUnlock_2[3:0] ? 1'h0 : _GEN_54; // @[elements.scala 190:33]
  wire  _GEN_71 = 4'h7 == idxUnlock_2[3:0] ? 1'h0 : _GEN_55; // @[elements.scala 190:33]
  wire  _GEN_72 = 4'h8 == idxUnlock_2[3:0] ? 1'h0 : _GEN_56; // @[elements.scala 190:33]
  wire  _GEN_73 = 4'h9 == idxUnlock_2[3:0] ? 1'h0 : _GEN_57; // @[elements.scala 190:33]
  wire  _GEN_74 = 4'ha == idxUnlock_2[3:0] ? 1'h0 : _GEN_58; // @[elements.scala 190:33]
  wire  _GEN_75 = 4'hb == idxUnlock_2[3:0] ? 1'h0 : _GEN_59; // @[elements.scala 190:33]
  wire  _GEN_76 = 4'hc == idxUnlock_2[3:0] ? 1'h0 : _GEN_60; // @[elements.scala 190:33]
  wire  _GEN_77 = 4'hd == idxUnlock_2[3:0] ? 1'h0 : _GEN_61; // @[elements.scala 190:33]
  wire  _GEN_78 = 4'he == idxUnlock_2[3:0] ? 1'h0 : _GEN_62; // @[elements.scala 190:33]
  wire  _GEN_79 = 4'hf == idxUnlock_2[3:0] ? 1'h0 : _GEN_63; // @[elements.scala 190:33]
  wire  _GEN_80 = _T_115 ? _GEN_64 : _GEN_48; // @[elements.scala 189:52]
  wire  _GEN_81 = _T_115 ? _GEN_65 : _GEN_49; // @[elements.scala 189:52]
  wire  _GEN_82 = _T_115 ? _GEN_66 : _GEN_50; // @[elements.scala 189:52]
  wire  _GEN_83 = _T_115 ? _GEN_67 : _GEN_51; // @[elements.scala 189:52]
  wire  _GEN_84 = _T_115 ? _GEN_68 : _GEN_52; // @[elements.scala 189:52]
  wire  _GEN_85 = _T_115 ? _GEN_69 : _GEN_53; // @[elements.scala 189:52]
  wire  _GEN_86 = _T_115 ? _GEN_70 : _GEN_54; // @[elements.scala 189:52]
  wire  _GEN_87 = _T_115 ? _GEN_71 : _GEN_55; // @[elements.scala 189:52]
  wire  _GEN_88 = _T_115 ? _GEN_72 : _GEN_56; // @[elements.scala 189:52]
  wire  _GEN_89 = _T_115 ? _GEN_73 : _GEN_57; // @[elements.scala 189:52]
  wire  _GEN_90 = _T_115 ? _GEN_74 : _GEN_58; // @[elements.scala 189:52]
  wire  _GEN_91 = _T_115 ? _GEN_75 : _GEN_59; // @[elements.scala 189:52]
  wire  _GEN_92 = _T_115 ? _GEN_76 : _GEN_60; // @[elements.scala 189:52]
  wire  _GEN_93 = _T_115 ? _GEN_77 : _GEN_61; // @[elements.scala 189:52]
  wire  _GEN_94 = _T_115 ? _GEN_78 : _GEN_62; // @[elements.scala 189:52]
  wire  _GEN_95 = _T_115 ? _GEN_79 : _GEN_63; // @[elements.scala 189:52]
  wire  _T_117 = io_unLock_3_in_valid & finder_3_io_value_valid; // @[elements.scala 189:23]
  wire [15:0] idxUnlock_3 = {{12'd0}, finder_3_io_value_bits}; // @[elements.scala 155:26 elements.scala 185:22]
  wire  _GEN_96 = 4'h0 == idxUnlock_3[3:0] ? 1'h0 : _GEN_80; // @[elements.scala 190:33]
  wire  _GEN_97 = 4'h1 == idxUnlock_3[3:0] ? 1'h0 : _GEN_81; // @[elements.scala 190:33]
  wire  _GEN_98 = 4'h2 == idxUnlock_3[3:0] ? 1'h0 : _GEN_82; // @[elements.scala 190:33]
  wire  _GEN_99 = 4'h3 == idxUnlock_3[3:0] ? 1'h0 : _GEN_83; // @[elements.scala 190:33]
  wire  _GEN_100 = 4'h4 == idxUnlock_3[3:0] ? 1'h0 : _GEN_84; // @[elements.scala 190:33]
  wire  _GEN_101 = 4'h5 == idxUnlock_3[3:0] ? 1'h0 : _GEN_85; // @[elements.scala 190:33]
  wire  _GEN_102 = 4'h6 == idxUnlock_3[3:0] ? 1'h0 : _GEN_86; // @[elements.scala 190:33]
  wire  _GEN_103 = 4'h7 == idxUnlock_3[3:0] ? 1'h0 : _GEN_87; // @[elements.scala 190:33]
  wire  _GEN_104 = 4'h8 == idxUnlock_3[3:0] ? 1'h0 : _GEN_88; // @[elements.scala 190:33]
  wire  _GEN_105 = 4'h9 == idxUnlock_3[3:0] ? 1'h0 : _GEN_89; // @[elements.scala 190:33]
  wire  _GEN_106 = 4'ha == idxUnlock_3[3:0] ? 1'h0 : _GEN_90; // @[elements.scala 190:33]
  wire  _GEN_107 = 4'hb == idxUnlock_3[3:0] ? 1'h0 : _GEN_91; // @[elements.scala 190:33]
  wire  _GEN_108 = 4'hc == idxUnlock_3[3:0] ? 1'h0 : _GEN_92; // @[elements.scala 190:33]
  wire  _GEN_109 = 4'hd == idxUnlock_3[3:0] ? 1'h0 : _GEN_93; // @[elements.scala 190:33]
  wire  _GEN_110 = 4'he == idxUnlock_3[3:0] ? 1'h0 : _GEN_94; // @[elements.scala 190:33]
  wire  _GEN_111 = 4'hf == idxUnlock_3[3:0] ? 1'h0 : _GEN_95; // @[elements.scala 190:33]
  wire  _GEN_112 = _T_117 ? _GEN_96 : _GEN_80; // @[elements.scala 189:52]
  wire  _GEN_113 = _T_117 ? _GEN_97 : _GEN_81; // @[elements.scala 189:52]
  wire  _GEN_114 = _T_117 ? _GEN_98 : _GEN_82; // @[elements.scala 189:52]
  wire  _GEN_115 = _T_117 ? _GEN_99 : _GEN_83; // @[elements.scala 189:52]
  wire  _GEN_116 = _T_117 ? _GEN_100 : _GEN_84; // @[elements.scala 189:52]
  wire  _GEN_117 = _T_117 ? _GEN_101 : _GEN_85; // @[elements.scala 189:52]
  wire  _GEN_118 = _T_117 ? _GEN_102 : _GEN_86; // @[elements.scala 189:52]
  wire  _GEN_119 = _T_117 ? _GEN_103 : _GEN_87; // @[elements.scala 189:52]
  wire  _GEN_120 = _T_117 ? _GEN_104 : _GEN_88; // @[elements.scala 189:52]
  wire  _GEN_121 = _T_117 ? _GEN_105 : _GEN_89; // @[elements.scala 189:52]
  wire  _GEN_122 = _T_117 ? _GEN_106 : _GEN_90; // @[elements.scala 189:52]
  wire  _GEN_123 = _T_117 ? _GEN_107 : _GEN_91; // @[elements.scala 189:52]
  wire  _GEN_124 = _T_117 ? _GEN_108 : _GEN_92; // @[elements.scala 189:52]
  wire  _GEN_125 = _T_117 ? _GEN_109 : _GEN_93; // @[elements.scala 189:52]
  wire  _GEN_126 = _T_117 ? _GEN_110 : _GEN_94; // @[elements.scala 189:52]
  wire  _GEN_127 = _T_117 ? _GEN_111 : _GEN_95; // @[elements.scala 189:52]
  wire  _T_119 = io_unLock_4_in_valid & finder_4_io_value_valid; // @[elements.scala 189:23]
  wire [15:0] idxUnlock_4 = {{12'd0}, finder_4_io_value_bits}; // @[elements.scala 155:26 elements.scala 185:22]
  wire  _GEN_128 = 4'h0 == idxUnlock_4[3:0] ? 1'h0 : _GEN_112; // @[elements.scala 190:33]
  wire  _GEN_129 = 4'h1 == idxUnlock_4[3:0] ? 1'h0 : _GEN_113; // @[elements.scala 190:33]
  wire  _GEN_130 = 4'h2 == idxUnlock_4[3:0] ? 1'h0 : _GEN_114; // @[elements.scala 190:33]
  wire  _GEN_131 = 4'h3 == idxUnlock_4[3:0] ? 1'h0 : _GEN_115; // @[elements.scala 190:33]
  wire  _GEN_132 = 4'h4 == idxUnlock_4[3:0] ? 1'h0 : _GEN_116; // @[elements.scala 190:33]
  wire  _GEN_133 = 4'h5 == idxUnlock_4[3:0] ? 1'h0 : _GEN_117; // @[elements.scala 190:33]
  wire  _GEN_134 = 4'h6 == idxUnlock_4[3:0] ? 1'h0 : _GEN_118; // @[elements.scala 190:33]
  wire  _GEN_135 = 4'h7 == idxUnlock_4[3:0] ? 1'h0 : _GEN_119; // @[elements.scala 190:33]
  wire  _GEN_136 = 4'h8 == idxUnlock_4[3:0] ? 1'h0 : _GEN_120; // @[elements.scala 190:33]
  wire  _GEN_137 = 4'h9 == idxUnlock_4[3:0] ? 1'h0 : _GEN_121; // @[elements.scala 190:33]
  wire  _GEN_138 = 4'ha == idxUnlock_4[3:0] ? 1'h0 : _GEN_122; // @[elements.scala 190:33]
  wire  _GEN_139 = 4'hb == idxUnlock_4[3:0] ? 1'h0 : _GEN_123; // @[elements.scala 190:33]
  wire  _GEN_140 = 4'hc == idxUnlock_4[3:0] ? 1'h0 : _GEN_124; // @[elements.scala 190:33]
  wire  _GEN_141 = 4'hd == idxUnlock_4[3:0] ? 1'h0 : _GEN_125; // @[elements.scala 190:33]
  wire  _GEN_142 = 4'he == idxUnlock_4[3:0] ? 1'h0 : _GEN_126; // @[elements.scala 190:33]
  wire  _GEN_143 = 4'hf == idxUnlock_4[3:0] ? 1'h0 : _GEN_127; // @[elements.scala 190:33]
  wire  _GEN_144 = _T_119 ? _GEN_128 : _GEN_112; // @[elements.scala 189:52]
  wire  _GEN_145 = _T_119 ? _GEN_129 : _GEN_113; // @[elements.scala 189:52]
  wire  _GEN_146 = _T_119 ? _GEN_130 : _GEN_114; // @[elements.scala 189:52]
  wire  _GEN_147 = _T_119 ? _GEN_131 : _GEN_115; // @[elements.scala 189:52]
  wire  _GEN_148 = _T_119 ? _GEN_132 : _GEN_116; // @[elements.scala 189:52]
  wire  _GEN_149 = _T_119 ? _GEN_133 : _GEN_117; // @[elements.scala 189:52]
  wire  _GEN_150 = _T_119 ? _GEN_134 : _GEN_118; // @[elements.scala 189:52]
  wire  _GEN_151 = _T_119 ? _GEN_135 : _GEN_119; // @[elements.scala 189:52]
  wire  _GEN_152 = _T_119 ? _GEN_136 : _GEN_120; // @[elements.scala 189:52]
  wire  _GEN_153 = _T_119 ? _GEN_137 : _GEN_121; // @[elements.scala 189:52]
  wire  _GEN_154 = _T_119 ? _GEN_138 : _GEN_122; // @[elements.scala 189:52]
  wire  _GEN_155 = _T_119 ? _GEN_139 : _GEN_123; // @[elements.scala 189:52]
  wire  _GEN_156 = _T_119 ? _GEN_140 : _GEN_124; // @[elements.scala 189:52]
  wire  _GEN_157 = _T_119 ? _GEN_141 : _GEN_125; // @[elements.scala 189:52]
  wire  _GEN_158 = _T_119 ? _GEN_142 : _GEN_126; // @[elements.scala 189:52]
  wire  _GEN_159 = _T_119 ? _GEN_143 : _GEN_127; // @[elements.scala 189:52]
  wire  _T_121 = io_unLock_5_in_valid & finder_5_io_value_valid; // @[elements.scala 189:23]
  wire [15:0] idxUnlock_5 = {{12'd0}, finder_5_io_value_bits}; // @[elements.scala 155:26 elements.scala 185:22]
  wire  _GEN_160 = 4'h0 == idxUnlock_5[3:0] ? 1'h0 : _GEN_144; // @[elements.scala 190:33]
  wire  _GEN_161 = 4'h1 == idxUnlock_5[3:0] ? 1'h0 : _GEN_145; // @[elements.scala 190:33]
  wire  _GEN_162 = 4'h2 == idxUnlock_5[3:0] ? 1'h0 : _GEN_146; // @[elements.scala 190:33]
  wire  _GEN_163 = 4'h3 == idxUnlock_5[3:0] ? 1'h0 : _GEN_147; // @[elements.scala 190:33]
  wire  _GEN_164 = 4'h4 == idxUnlock_5[3:0] ? 1'h0 : _GEN_148; // @[elements.scala 190:33]
  wire  _GEN_165 = 4'h5 == idxUnlock_5[3:0] ? 1'h0 : _GEN_149; // @[elements.scala 190:33]
  wire  _GEN_166 = 4'h6 == idxUnlock_5[3:0] ? 1'h0 : _GEN_150; // @[elements.scala 190:33]
  wire  _GEN_167 = 4'h7 == idxUnlock_5[3:0] ? 1'h0 : _GEN_151; // @[elements.scala 190:33]
  wire  _GEN_168 = 4'h8 == idxUnlock_5[3:0] ? 1'h0 : _GEN_152; // @[elements.scala 190:33]
  wire  _GEN_169 = 4'h9 == idxUnlock_5[3:0] ? 1'h0 : _GEN_153; // @[elements.scala 190:33]
  wire  _GEN_170 = 4'ha == idxUnlock_5[3:0] ? 1'h0 : _GEN_154; // @[elements.scala 190:33]
  wire  _GEN_171 = 4'hb == idxUnlock_5[3:0] ? 1'h0 : _GEN_155; // @[elements.scala 190:33]
  wire  _GEN_172 = 4'hc == idxUnlock_5[3:0] ? 1'h0 : _GEN_156; // @[elements.scala 190:33]
  wire  _GEN_173 = 4'hd == idxUnlock_5[3:0] ? 1'h0 : _GEN_157; // @[elements.scala 190:33]
  wire  _GEN_174 = 4'he == idxUnlock_5[3:0] ? 1'h0 : _GEN_158; // @[elements.scala 190:33]
  wire  _GEN_175 = 4'hf == idxUnlock_5[3:0] ? 1'h0 : _GEN_159; // @[elements.scala 190:33]
  wire  _GEN_176 = _T_121 ? _GEN_160 : _GEN_144; // @[elements.scala 189:52]
  wire  _GEN_177 = _T_121 ? _GEN_161 : _GEN_145; // @[elements.scala 189:52]
  wire  _GEN_178 = _T_121 ? _GEN_162 : _GEN_146; // @[elements.scala 189:52]
  wire  _GEN_179 = _T_121 ? _GEN_163 : _GEN_147; // @[elements.scala 189:52]
  wire  _GEN_180 = _T_121 ? _GEN_164 : _GEN_148; // @[elements.scala 189:52]
  wire  _GEN_181 = _T_121 ? _GEN_165 : _GEN_149; // @[elements.scala 189:52]
  wire  _GEN_182 = _T_121 ? _GEN_166 : _GEN_150; // @[elements.scala 189:52]
  wire  _GEN_183 = _T_121 ? _GEN_167 : _GEN_151; // @[elements.scala 189:52]
  wire  _GEN_184 = _T_121 ? _GEN_168 : _GEN_152; // @[elements.scala 189:52]
  wire  _GEN_185 = _T_121 ? _GEN_169 : _GEN_153; // @[elements.scala 189:52]
  wire  _GEN_186 = _T_121 ? _GEN_170 : _GEN_154; // @[elements.scala 189:52]
  wire  _GEN_187 = _T_121 ? _GEN_171 : _GEN_155; // @[elements.scala 189:52]
  wire  _GEN_188 = _T_121 ? _GEN_172 : _GEN_156; // @[elements.scala 189:52]
  wire  _GEN_189 = _T_121 ? _GEN_173 : _GEN_157; // @[elements.scala 189:52]
  wire  _GEN_190 = _T_121 ? _GEN_174 : _GEN_158; // @[elements.scala 189:52]
  wire  _GEN_191 = _T_121 ? _GEN_175 : _GEN_159; // @[elements.scala 189:52]
  wire  _T_123 = io_unLock_6_in_valid & finder_6_io_value_valid; // @[elements.scala 189:23]
  wire [15:0] idxUnlock_6 = {{12'd0}, finder_6_io_value_bits}; // @[elements.scala 155:26 elements.scala 185:22]
  wire  _GEN_192 = 4'h0 == idxUnlock_6[3:0] ? 1'h0 : _GEN_176; // @[elements.scala 190:33]
  wire  _GEN_193 = 4'h1 == idxUnlock_6[3:0] ? 1'h0 : _GEN_177; // @[elements.scala 190:33]
  wire  _GEN_194 = 4'h2 == idxUnlock_6[3:0] ? 1'h0 : _GEN_178; // @[elements.scala 190:33]
  wire  _GEN_195 = 4'h3 == idxUnlock_6[3:0] ? 1'h0 : _GEN_179; // @[elements.scala 190:33]
  wire  _GEN_196 = 4'h4 == idxUnlock_6[3:0] ? 1'h0 : _GEN_180; // @[elements.scala 190:33]
  wire  _GEN_197 = 4'h5 == idxUnlock_6[3:0] ? 1'h0 : _GEN_181; // @[elements.scala 190:33]
  wire  _GEN_198 = 4'h6 == idxUnlock_6[3:0] ? 1'h0 : _GEN_182; // @[elements.scala 190:33]
  wire  _GEN_199 = 4'h7 == idxUnlock_6[3:0] ? 1'h0 : _GEN_183; // @[elements.scala 190:33]
  wire  _GEN_200 = 4'h8 == idxUnlock_6[3:0] ? 1'h0 : _GEN_184; // @[elements.scala 190:33]
  wire  _GEN_201 = 4'h9 == idxUnlock_6[3:0] ? 1'h0 : _GEN_185; // @[elements.scala 190:33]
  wire  _GEN_202 = 4'ha == idxUnlock_6[3:0] ? 1'h0 : _GEN_186; // @[elements.scala 190:33]
  wire  _GEN_203 = 4'hb == idxUnlock_6[3:0] ? 1'h0 : _GEN_187; // @[elements.scala 190:33]
  wire  _GEN_204 = 4'hc == idxUnlock_6[3:0] ? 1'h0 : _GEN_188; // @[elements.scala 190:33]
  wire  _GEN_205 = 4'hd == idxUnlock_6[3:0] ? 1'h0 : _GEN_189; // @[elements.scala 190:33]
  wire  _GEN_206 = 4'he == idxUnlock_6[3:0] ? 1'h0 : _GEN_190; // @[elements.scala 190:33]
  wire  _GEN_207 = 4'hf == idxUnlock_6[3:0] ? 1'h0 : _GEN_191; // @[elements.scala 190:33]
  wire  _GEN_208 = _T_123 ? _GEN_192 : _GEN_176; // @[elements.scala 189:52]
  wire  _GEN_209 = _T_123 ? _GEN_193 : _GEN_177; // @[elements.scala 189:52]
  wire  _GEN_210 = _T_123 ? _GEN_194 : _GEN_178; // @[elements.scala 189:52]
  wire  _GEN_211 = _T_123 ? _GEN_195 : _GEN_179; // @[elements.scala 189:52]
  wire  _GEN_212 = _T_123 ? _GEN_196 : _GEN_180; // @[elements.scala 189:52]
  wire  _GEN_213 = _T_123 ? _GEN_197 : _GEN_181; // @[elements.scala 189:52]
  wire  _GEN_214 = _T_123 ? _GEN_198 : _GEN_182; // @[elements.scala 189:52]
  wire  _GEN_215 = _T_123 ? _GEN_199 : _GEN_183; // @[elements.scala 189:52]
  wire  _GEN_216 = _T_123 ? _GEN_200 : _GEN_184; // @[elements.scala 189:52]
  wire  _GEN_217 = _T_123 ? _GEN_201 : _GEN_185; // @[elements.scala 189:52]
  wire  _GEN_218 = _T_123 ? _GEN_202 : _GEN_186; // @[elements.scala 189:52]
  wire  _GEN_219 = _T_123 ? _GEN_203 : _GEN_187; // @[elements.scala 189:52]
  wire  _GEN_220 = _T_123 ? _GEN_204 : _GEN_188; // @[elements.scala 189:52]
  wire  _GEN_221 = _T_123 ? _GEN_205 : _GEN_189; // @[elements.scala 189:52]
  wire  _GEN_222 = _T_123 ? _GEN_206 : _GEN_190; // @[elements.scala 189:52]
  wire  _GEN_223 = _T_123 ? _GEN_207 : _GEN_191; // @[elements.scala 189:52]
  wire  _T_125 = io_unLock_7_in_valid & finder_7_io_value_valid; // @[elements.scala 189:23]
  wire [15:0] idxUnlock_7 = {{12'd0}, finder_7_io_value_bits}; // @[elements.scala 155:26 elements.scala 185:22]
  wire  _GEN_224 = 4'h0 == idxUnlock_7[3:0] ? 1'h0 : _GEN_208; // @[elements.scala 190:33]
  wire  _GEN_225 = 4'h1 == idxUnlock_7[3:0] ? 1'h0 : _GEN_209; // @[elements.scala 190:33]
  wire  _GEN_226 = 4'h2 == idxUnlock_7[3:0] ? 1'h0 : _GEN_210; // @[elements.scala 190:33]
  wire  _GEN_227 = 4'h3 == idxUnlock_7[3:0] ? 1'h0 : _GEN_211; // @[elements.scala 190:33]
  wire  _GEN_228 = 4'h4 == idxUnlock_7[3:0] ? 1'h0 : _GEN_212; // @[elements.scala 190:33]
  wire  _GEN_229 = 4'h5 == idxUnlock_7[3:0] ? 1'h0 : _GEN_213; // @[elements.scala 190:33]
  wire  _GEN_230 = 4'h6 == idxUnlock_7[3:0] ? 1'h0 : _GEN_214; // @[elements.scala 190:33]
  wire  _GEN_231 = 4'h7 == idxUnlock_7[3:0] ? 1'h0 : _GEN_215; // @[elements.scala 190:33]
  wire  _GEN_232 = 4'h8 == idxUnlock_7[3:0] ? 1'h0 : _GEN_216; // @[elements.scala 190:33]
  wire  _GEN_233 = 4'h9 == idxUnlock_7[3:0] ? 1'h0 : _GEN_217; // @[elements.scala 190:33]
  wire  _GEN_234 = 4'ha == idxUnlock_7[3:0] ? 1'h0 : _GEN_218; // @[elements.scala 190:33]
  wire  _GEN_235 = 4'hb == idxUnlock_7[3:0] ? 1'h0 : _GEN_219; // @[elements.scala 190:33]
  wire  _GEN_236 = 4'hc == idxUnlock_7[3:0] ? 1'h0 : _GEN_220; // @[elements.scala 190:33]
  wire  _GEN_237 = 4'hd == idxUnlock_7[3:0] ? 1'h0 : _GEN_221; // @[elements.scala 190:33]
  wire  _GEN_238 = 4'he == idxUnlock_7[3:0] ? 1'h0 : _GEN_222; // @[elements.scala 190:33]
  wire  _GEN_239 = 4'hf == idxUnlock_7[3:0] ? 1'h0 : _GEN_223; // @[elements.scala 190:33]
  wire  _GEN_240 = _T_125 ? _GEN_224 : _GEN_208; // @[elements.scala 189:52]
  wire  _GEN_241 = _T_125 ? _GEN_225 : _GEN_209; // @[elements.scala 189:52]
  wire  _GEN_242 = _T_125 ? _GEN_226 : _GEN_210; // @[elements.scala 189:52]
  wire  _GEN_243 = _T_125 ? _GEN_227 : _GEN_211; // @[elements.scala 189:52]
  wire  _GEN_244 = _T_125 ? _GEN_228 : _GEN_212; // @[elements.scala 189:52]
  wire  _GEN_245 = _T_125 ? _GEN_229 : _GEN_213; // @[elements.scala 189:52]
  wire  _GEN_246 = _T_125 ? _GEN_230 : _GEN_214; // @[elements.scala 189:52]
  wire  _GEN_247 = _T_125 ? _GEN_231 : _GEN_215; // @[elements.scala 189:52]
  wire  _GEN_248 = _T_125 ? _GEN_232 : _GEN_216; // @[elements.scala 189:52]
  wire  _GEN_249 = _T_125 ? _GEN_233 : _GEN_217; // @[elements.scala 189:52]
  wire  _GEN_250 = _T_125 ? _GEN_234 : _GEN_218; // @[elements.scala 189:52]
  wire  _GEN_251 = _T_125 ? _GEN_235 : _GEN_219; // @[elements.scala 189:52]
  wire  _GEN_252 = _T_125 ? _GEN_236 : _GEN_220; // @[elements.scala 189:52]
  wire  _GEN_253 = _T_125 ? _GEN_237 : _GEN_221; // @[elements.scala 189:52]
  wire  _GEN_254 = _T_125 ? _GEN_238 : _GEN_222; // @[elements.scala 189:52]
  wire  _GEN_255 = _T_125 ? _GEN_239 : _GEN_223; // @[elements.scala 189:52]
  wire  _T_127 = ~valid_0; // @[elements.scala 196:46]
  wire  _T_128 = ~valid_1; // @[elements.scala 196:46]
  wire  _T_129 = ~valid_2; // @[elements.scala 196:46]
  wire  _T_130 = ~valid_3; // @[elements.scala 196:46]
  wire  _T_131 = ~valid_4; // @[elements.scala 196:46]
  wire  _T_132 = ~valid_5; // @[elements.scala 196:46]
  wire  _T_133 = ~valid_6; // @[elements.scala 196:46]
  wire  _T_134 = ~valid_7; // @[elements.scala 196:46]
  wire  _T_135 = ~valid_8; // @[elements.scala 196:46]
  wire  _T_136 = ~valid_9; // @[elements.scala 196:46]
  wire  _T_137 = ~valid_10; // @[elements.scala 196:46]
  wire  _T_138 = ~valid_11; // @[elements.scala 196:46]
  wire  _T_139 = ~valid_12; // @[elements.scala 196:46]
  wire  _T_140 = ~valid_13; // @[elements.scala 196:46]
  wire  _T_141 = ~valid_14; // @[elements.scala 196:46]
  wire  _T_142 = ~valid_15; // @[elements.scala 196:46]
  wire [4:0] _GEN_256 = _T_142 ? 5'hf : 5'h10; // @[elements.scala 196:59]
  wire [4:0] _GEN_257 = _T_141 ? 5'he : _GEN_256; // @[elements.scala 196:59]
  wire [4:0] _GEN_258 = _T_140 ? 5'hd : _GEN_257; // @[elements.scala 196:59]
  wire [4:0] _GEN_259 = _T_139 ? 5'hc : _GEN_258; // @[elements.scala 196:59]
  wire [4:0] _GEN_260 = _T_138 ? 5'hb : _GEN_259; // @[elements.scala 196:59]
  wire [4:0] _GEN_261 = _T_137 ? 5'ha : _GEN_260; // @[elements.scala 196:59]
  wire [4:0] _GEN_262 = _T_136 ? 5'h9 : _GEN_261; // @[elements.scala 196:59]
  wire [4:0] _GEN_263 = _T_135 ? 5'h8 : _GEN_262; // @[elements.scala 196:59]
  wire [4:0] _GEN_264 = _T_134 ? 5'h7 : _GEN_263; // @[elements.scala 196:59]
  wire [4:0] _GEN_265 = _T_133 ? 5'h6 : _GEN_264; // @[elements.scala 196:59]
  wire [4:0] _GEN_266 = _T_132 ? 5'h5 : _GEN_265; // @[elements.scala 196:59]
  wire [4:0] _GEN_267 = _T_131 ? 5'h4 : _GEN_266; // @[elements.scala 196:59]
  wire [4:0] _GEN_268 = _T_130 ? 5'h3 : _GEN_267; // @[elements.scala 196:59]
  wire [4:0] _GEN_269 = _T_129 ? 5'h2 : _GEN_268; // @[elements.scala 196:59]
  wire [4:0] _GEN_270 = _T_128 ? 5'h1 : _GEN_269; // @[elements.scala 196:59]
  wire [4:0] _GEN_271 = _T_127 ? 5'h0 : _GEN_270; // @[elements.scala 196:59]
  wire [15:0] idxLocking = {{11'd0}, _GEN_271}; // @[elements.scala 153:26 elements.scala 177:16 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28]
  wire  _GEN_337 = 4'h0 == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_305 = _GEN_337 | _GEN_240; // @[elements.scala 212:27]
  wire  _GEN_338 = 4'h1 == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_306 = _GEN_338 | _GEN_241; // @[elements.scala 212:27]
  wire  _GEN_339 = 4'h2 == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_307 = _GEN_339 | _GEN_242; // @[elements.scala 212:27]
  wire  _GEN_340 = 4'h3 == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_308 = _GEN_340 | _GEN_243; // @[elements.scala 212:27]
  wire  _GEN_341 = 4'h4 == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_309 = _GEN_341 | _GEN_244; // @[elements.scala 212:27]
  wire  _GEN_342 = 4'h5 == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_310 = _GEN_342 | _GEN_245; // @[elements.scala 212:27]
  wire  _GEN_343 = 4'h6 == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_311 = _GEN_343 | _GEN_246; // @[elements.scala 212:27]
  wire  _GEN_344 = 4'h7 == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_312 = _GEN_344 | _GEN_247; // @[elements.scala 212:27]
  wire  _GEN_345 = 4'h8 == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_313 = _GEN_345 | _GEN_248; // @[elements.scala 212:27]
  wire  _GEN_346 = 4'h9 == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_314 = _GEN_346 | _GEN_249; // @[elements.scala 212:27]
  wire  _GEN_347 = 4'ha == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_315 = _GEN_347 | _GEN_250; // @[elements.scala 212:27]
  wire  _GEN_348 = 4'hb == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_316 = _GEN_348 | _GEN_251; // @[elements.scala 212:27]
  wire  _GEN_349 = 4'hc == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_317 = _GEN_349 | _GEN_252; // @[elements.scala 212:27]
  wire  _GEN_350 = 4'hd == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_318 = _GEN_350 | _GEN_253; // @[elements.scala 212:27]
  wire  _GEN_351 = 4'he == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_319 = _GEN_351 | _GEN_254; // @[elements.scala 212:27]
  wire  _GEN_352 = 4'hf == idxLocking[3:0]; // @[elements.scala 212:27]
  wire  _GEN_320 = _GEN_352 | _GEN_255; // @[elements.scala 212:27]
  Find_9 finder_0 ( // @[elements.scala 158:28]
    .io_key(finder_0_io_key),
    .io_data_0(finder_0_io_data_0),
    .io_data_1(finder_0_io_data_1),
    .io_data_2(finder_0_io_data_2),
    .io_data_3(finder_0_io_data_3),
    .io_data_4(finder_0_io_data_4),
    .io_data_5(finder_0_io_data_5),
    .io_data_6(finder_0_io_data_6),
    .io_data_7(finder_0_io_data_7),
    .io_data_8(finder_0_io_data_8),
    .io_data_9(finder_0_io_data_9),
    .io_data_10(finder_0_io_data_10),
    .io_data_11(finder_0_io_data_11),
    .io_data_12(finder_0_io_data_12),
    .io_data_13(finder_0_io_data_13),
    .io_data_14(finder_0_io_data_14),
    .io_data_15(finder_0_io_data_15),
    .io_valid_0(finder_0_io_valid_0),
    .io_valid_1(finder_0_io_valid_1),
    .io_valid_2(finder_0_io_valid_2),
    .io_valid_3(finder_0_io_valid_3),
    .io_valid_4(finder_0_io_valid_4),
    .io_valid_5(finder_0_io_valid_5),
    .io_valid_6(finder_0_io_valid_6),
    .io_valid_7(finder_0_io_valid_7),
    .io_valid_8(finder_0_io_valid_8),
    .io_valid_9(finder_0_io_valid_9),
    .io_valid_10(finder_0_io_valid_10),
    .io_valid_11(finder_0_io_valid_11),
    .io_valid_12(finder_0_io_valid_12),
    .io_valid_13(finder_0_io_valid_13),
    .io_valid_14(finder_0_io_valid_14),
    .io_valid_15(finder_0_io_valid_15),
    .io_value_valid(finder_0_io_value_valid),
    .io_value_bits(finder_0_io_value_bits)
  );
  Find_9 finder_1 ( // @[elements.scala 158:28]
    .io_key(finder_1_io_key),
    .io_data_0(finder_1_io_data_0),
    .io_data_1(finder_1_io_data_1),
    .io_data_2(finder_1_io_data_2),
    .io_data_3(finder_1_io_data_3),
    .io_data_4(finder_1_io_data_4),
    .io_data_5(finder_1_io_data_5),
    .io_data_6(finder_1_io_data_6),
    .io_data_7(finder_1_io_data_7),
    .io_data_8(finder_1_io_data_8),
    .io_data_9(finder_1_io_data_9),
    .io_data_10(finder_1_io_data_10),
    .io_data_11(finder_1_io_data_11),
    .io_data_12(finder_1_io_data_12),
    .io_data_13(finder_1_io_data_13),
    .io_data_14(finder_1_io_data_14),
    .io_data_15(finder_1_io_data_15),
    .io_valid_0(finder_1_io_valid_0),
    .io_valid_1(finder_1_io_valid_1),
    .io_valid_2(finder_1_io_valid_2),
    .io_valid_3(finder_1_io_valid_3),
    .io_valid_4(finder_1_io_valid_4),
    .io_valid_5(finder_1_io_valid_5),
    .io_valid_6(finder_1_io_valid_6),
    .io_valid_7(finder_1_io_valid_7),
    .io_valid_8(finder_1_io_valid_8),
    .io_valid_9(finder_1_io_valid_9),
    .io_valid_10(finder_1_io_valid_10),
    .io_valid_11(finder_1_io_valid_11),
    .io_valid_12(finder_1_io_valid_12),
    .io_valid_13(finder_1_io_valid_13),
    .io_valid_14(finder_1_io_valid_14),
    .io_valid_15(finder_1_io_valid_15),
    .io_value_valid(finder_1_io_value_valid),
    .io_value_bits(finder_1_io_value_bits)
  );
  Find_9 finder_2 ( // @[elements.scala 158:28]
    .io_key(finder_2_io_key),
    .io_data_0(finder_2_io_data_0),
    .io_data_1(finder_2_io_data_1),
    .io_data_2(finder_2_io_data_2),
    .io_data_3(finder_2_io_data_3),
    .io_data_4(finder_2_io_data_4),
    .io_data_5(finder_2_io_data_5),
    .io_data_6(finder_2_io_data_6),
    .io_data_7(finder_2_io_data_7),
    .io_data_8(finder_2_io_data_8),
    .io_data_9(finder_2_io_data_9),
    .io_data_10(finder_2_io_data_10),
    .io_data_11(finder_2_io_data_11),
    .io_data_12(finder_2_io_data_12),
    .io_data_13(finder_2_io_data_13),
    .io_data_14(finder_2_io_data_14),
    .io_data_15(finder_2_io_data_15),
    .io_valid_0(finder_2_io_valid_0),
    .io_valid_1(finder_2_io_valid_1),
    .io_valid_2(finder_2_io_valid_2),
    .io_valid_3(finder_2_io_valid_3),
    .io_valid_4(finder_2_io_valid_4),
    .io_valid_5(finder_2_io_valid_5),
    .io_valid_6(finder_2_io_valid_6),
    .io_valid_7(finder_2_io_valid_7),
    .io_valid_8(finder_2_io_valid_8),
    .io_valid_9(finder_2_io_valid_9),
    .io_valid_10(finder_2_io_valid_10),
    .io_valid_11(finder_2_io_valid_11),
    .io_valid_12(finder_2_io_valid_12),
    .io_valid_13(finder_2_io_valid_13),
    .io_valid_14(finder_2_io_valid_14),
    .io_valid_15(finder_2_io_valid_15),
    .io_value_valid(finder_2_io_value_valid),
    .io_value_bits(finder_2_io_value_bits)
  );
  Find_9 finder_3 ( // @[elements.scala 158:28]
    .io_key(finder_3_io_key),
    .io_data_0(finder_3_io_data_0),
    .io_data_1(finder_3_io_data_1),
    .io_data_2(finder_3_io_data_2),
    .io_data_3(finder_3_io_data_3),
    .io_data_4(finder_3_io_data_4),
    .io_data_5(finder_3_io_data_5),
    .io_data_6(finder_3_io_data_6),
    .io_data_7(finder_3_io_data_7),
    .io_data_8(finder_3_io_data_8),
    .io_data_9(finder_3_io_data_9),
    .io_data_10(finder_3_io_data_10),
    .io_data_11(finder_3_io_data_11),
    .io_data_12(finder_3_io_data_12),
    .io_data_13(finder_3_io_data_13),
    .io_data_14(finder_3_io_data_14),
    .io_data_15(finder_3_io_data_15),
    .io_valid_0(finder_3_io_valid_0),
    .io_valid_1(finder_3_io_valid_1),
    .io_valid_2(finder_3_io_valid_2),
    .io_valid_3(finder_3_io_valid_3),
    .io_valid_4(finder_3_io_valid_4),
    .io_valid_5(finder_3_io_valid_5),
    .io_valid_6(finder_3_io_valid_6),
    .io_valid_7(finder_3_io_valid_7),
    .io_valid_8(finder_3_io_valid_8),
    .io_valid_9(finder_3_io_valid_9),
    .io_valid_10(finder_3_io_valid_10),
    .io_valid_11(finder_3_io_valid_11),
    .io_valid_12(finder_3_io_valid_12),
    .io_valid_13(finder_3_io_valid_13),
    .io_valid_14(finder_3_io_valid_14),
    .io_valid_15(finder_3_io_valid_15),
    .io_value_valid(finder_3_io_value_valid),
    .io_value_bits(finder_3_io_value_bits)
  );
  Find_9 finder_4 ( // @[elements.scala 158:28]
    .io_key(finder_4_io_key),
    .io_data_0(finder_4_io_data_0),
    .io_data_1(finder_4_io_data_1),
    .io_data_2(finder_4_io_data_2),
    .io_data_3(finder_4_io_data_3),
    .io_data_4(finder_4_io_data_4),
    .io_data_5(finder_4_io_data_5),
    .io_data_6(finder_4_io_data_6),
    .io_data_7(finder_4_io_data_7),
    .io_data_8(finder_4_io_data_8),
    .io_data_9(finder_4_io_data_9),
    .io_data_10(finder_4_io_data_10),
    .io_data_11(finder_4_io_data_11),
    .io_data_12(finder_4_io_data_12),
    .io_data_13(finder_4_io_data_13),
    .io_data_14(finder_4_io_data_14),
    .io_data_15(finder_4_io_data_15),
    .io_valid_0(finder_4_io_valid_0),
    .io_valid_1(finder_4_io_valid_1),
    .io_valid_2(finder_4_io_valid_2),
    .io_valid_3(finder_4_io_valid_3),
    .io_valid_4(finder_4_io_valid_4),
    .io_valid_5(finder_4_io_valid_5),
    .io_valid_6(finder_4_io_valid_6),
    .io_valid_7(finder_4_io_valid_7),
    .io_valid_8(finder_4_io_valid_8),
    .io_valid_9(finder_4_io_valid_9),
    .io_valid_10(finder_4_io_valid_10),
    .io_valid_11(finder_4_io_valid_11),
    .io_valid_12(finder_4_io_valid_12),
    .io_valid_13(finder_4_io_valid_13),
    .io_valid_14(finder_4_io_valid_14),
    .io_valid_15(finder_4_io_valid_15),
    .io_value_valid(finder_4_io_value_valid),
    .io_value_bits(finder_4_io_value_bits)
  );
  Find_9 finder_5 ( // @[elements.scala 158:28]
    .io_key(finder_5_io_key),
    .io_data_0(finder_5_io_data_0),
    .io_data_1(finder_5_io_data_1),
    .io_data_2(finder_5_io_data_2),
    .io_data_3(finder_5_io_data_3),
    .io_data_4(finder_5_io_data_4),
    .io_data_5(finder_5_io_data_5),
    .io_data_6(finder_5_io_data_6),
    .io_data_7(finder_5_io_data_7),
    .io_data_8(finder_5_io_data_8),
    .io_data_9(finder_5_io_data_9),
    .io_data_10(finder_5_io_data_10),
    .io_data_11(finder_5_io_data_11),
    .io_data_12(finder_5_io_data_12),
    .io_data_13(finder_5_io_data_13),
    .io_data_14(finder_5_io_data_14),
    .io_data_15(finder_5_io_data_15),
    .io_valid_0(finder_5_io_valid_0),
    .io_valid_1(finder_5_io_valid_1),
    .io_valid_2(finder_5_io_valid_2),
    .io_valid_3(finder_5_io_valid_3),
    .io_valid_4(finder_5_io_valid_4),
    .io_valid_5(finder_5_io_valid_5),
    .io_valid_6(finder_5_io_valid_6),
    .io_valid_7(finder_5_io_valid_7),
    .io_valid_8(finder_5_io_valid_8),
    .io_valid_9(finder_5_io_valid_9),
    .io_valid_10(finder_5_io_valid_10),
    .io_valid_11(finder_5_io_valid_11),
    .io_valid_12(finder_5_io_valid_12),
    .io_valid_13(finder_5_io_valid_13),
    .io_valid_14(finder_5_io_valid_14),
    .io_valid_15(finder_5_io_valid_15),
    .io_value_valid(finder_5_io_value_valid),
    .io_value_bits(finder_5_io_value_bits)
  );
  Find_9 finder_6 ( // @[elements.scala 158:28]
    .io_key(finder_6_io_key),
    .io_data_0(finder_6_io_data_0),
    .io_data_1(finder_6_io_data_1),
    .io_data_2(finder_6_io_data_2),
    .io_data_3(finder_6_io_data_3),
    .io_data_4(finder_6_io_data_4),
    .io_data_5(finder_6_io_data_5),
    .io_data_6(finder_6_io_data_6),
    .io_data_7(finder_6_io_data_7),
    .io_data_8(finder_6_io_data_8),
    .io_data_9(finder_6_io_data_9),
    .io_data_10(finder_6_io_data_10),
    .io_data_11(finder_6_io_data_11),
    .io_data_12(finder_6_io_data_12),
    .io_data_13(finder_6_io_data_13),
    .io_data_14(finder_6_io_data_14),
    .io_data_15(finder_6_io_data_15),
    .io_valid_0(finder_6_io_valid_0),
    .io_valid_1(finder_6_io_valid_1),
    .io_valid_2(finder_6_io_valid_2),
    .io_valid_3(finder_6_io_valid_3),
    .io_valid_4(finder_6_io_valid_4),
    .io_valid_5(finder_6_io_valid_5),
    .io_valid_6(finder_6_io_valid_6),
    .io_valid_7(finder_6_io_valid_7),
    .io_valid_8(finder_6_io_valid_8),
    .io_valid_9(finder_6_io_valid_9),
    .io_valid_10(finder_6_io_valid_10),
    .io_valid_11(finder_6_io_valid_11),
    .io_valid_12(finder_6_io_valid_12),
    .io_valid_13(finder_6_io_valid_13),
    .io_valid_14(finder_6_io_valid_14),
    .io_valid_15(finder_6_io_valid_15),
    .io_value_valid(finder_6_io_value_valid),
    .io_value_bits(finder_6_io_value_bits)
  );
  Find_9 finder_7 ( // @[elements.scala 158:28]
    .io_key(finder_7_io_key),
    .io_data_0(finder_7_io_data_0),
    .io_data_1(finder_7_io_data_1),
    .io_data_2(finder_7_io_data_2),
    .io_data_3(finder_7_io_data_3),
    .io_data_4(finder_7_io_data_4),
    .io_data_5(finder_7_io_data_5),
    .io_data_6(finder_7_io_data_6),
    .io_data_7(finder_7_io_data_7),
    .io_data_8(finder_7_io_data_8),
    .io_data_9(finder_7_io_data_9),
    .io_data_10(finder_7_io_data_10),
    .io_data_11(finder_7_io_data_11),
    .io_data_12(finder_7_io_data_12),
    .io_data_13(finder_7_io_data_13),
    .io_data_14(finder_7_io_data_14),
    .io_data_15(finder_7_io_data_15),
    .io_valid_0(finder_7_io_valid_0),
    .io_valid_1(finder_7_io_valid_1),
    .io_valid_2(finder_7_io_valid_2),
    .io_valid_3(finder_7_io_valid_3),
    .io_valid_4(finder_7_io_valid_4),
    .io_valid_5(finder_7_io_valid_5),
    .io_valid_6(finder_7_io_valid_6),
    .io_valid_7(finder_7_io_valid_7),
    .io_valid_8(finder_7_io_valid_8),
    .io_valid_9(finder_7_io_valid_9),
    .io_valid_10(finder_7_io_valid_10),
    .io_valid_11(finder_7_io_valid_11),
    .io_valid_12(finder_7_io_valid_12),
    .io_valid_13(finder_7_io_valid_13),
    .io_valid_14(finder_7_io_valid_14),
    .io_valid_15(finder_7_io_valid_15),
    .io_value_valid(finder_7_io_value_valid),
    .io_value_bits(finder_7_io_value_bits)
  );
  assign io_probe_out_valid = io_probe_in_valid; // @[elements.scala 203:24]
  assign io_probe_out_bits = _T_158 != 16'h0; // @[elements.scala 202:23]
  assign finder_0_io_key = io_unLock_0_in_bits_addr; // @[elements.scala 183:26]
  assign finder_0_io_data_0 = addrVec_0; // @[elements.scala 182:27]
  assign finder_0_io_data_1 = addrVec_1; // @[elements.scala 182:27]
  assign finder_0_io_data_2 = addrVec_2; // @[elements.scala 182:27]
  assign finder_0_io_data_3 = addrVec_3; // @[elements.scala 182:27]
  assign finder_0_io_data_4 = addrVec_4; // @[elements.scala 182:27]
  assign finder_0_io_data_5 = addrVec_5; // @[elements.scala 182:27]
  assign finder_0_io_data_6 = addrVec_6; // @[elements.scala 182:27]
  assign finder_0_io_data_7 = addrVec_7; // @[elements.scala 182:27]
  assign finder_0_io_data_8 = addrVec_8; // @[elements.scala 182:27]
  assign finder_0_io_data_9 = addrVec_9; // @[elements.scala 182:27]
  assign finder_0_io_data_10 = addrVec_10; // @[elements.scala 182:27]
  assign finder_0_io_data_11 = addrVec_11; // @[elements.scala 182:27]
  assign finder_0_io_data_12 = addrVec_12; // @[elements.scala 182:27]
  assign finder_0_io_data_13 = addrVec_13; // @[elements.scala 182:27]
  assign finder_0_io_data_14 = addrVec_14; // @[elements.scala 182:27]
  assign finder_0_io_data_15 = addrVec_15; // @[elements.scala 182:27]
  assign finder_0_io_valid_0 = valid_0; // @[elements.scala 184:28]
  assign finder_0_io_valid_1 = valid_1; // @[elements.scala 184:28]
  assign finder_0_io_valid_2 = valid_2; // @[elements.scala 184:28]
  assign finder_0_io_valid_3 = valid_3; // @[elements.scala 184:28]
  assign finder_0_io_valid_4 = valid_4; // @[elements.scala 184:28]
  assign finder_0_io_valid_5 = valid_5; // @[elements.scala 184:28]
  assign finder_0_io_valid_6 = valid_6; // @[elements.scala 184:28]
  assign finder_0_io_valid_7 = valid_7; // @[elements.scala 184:28]
  assign finder_0_io_valid_8 = valid_8; // @[elements.scala 184:28]
  assign finder_0_io_valid_9 = valid_9; // @[elements.scala 184:28]
  assign finder_0_io_valid_10 = valid_10; // @[elements.scala 184:28]
  assign finder_0_io_valid_11 = valid_11; // @[elements.scala 184:28]
  assign finder_0_io_valid_12 = valid_12; // @[elements.scala 184:28]
  assign finder_0_io_valid_13 = valid_13; // @[elements.scala 184:28]
  assign finder_0_io_valid_14 = valid_14; // @[elements.scala 184:28]
  assign finder_0_io_valid_15 = valid_15; // @[elements.scala 184:28]
  assign finder_1_io_key = io_unLock_1_in_bits_addr; // @[elements.scala 183:26]
  assign finder_1_io_data_0 = addrVec_0; // @[elements.scala 182:27]
  assign finder_1_io_data_1 = addrVec_1; // @[elements.scala 182:27]
  assign finder_1_io_data_2 = addrVec_2; // @[elements.scala 182:27]
  assign finder_1_io_data_3 = addrVec_3; // @[elements.scala 182:27]
  assign finder_1_io_data_4 = addrVec_4; // @[elements.scala 182:27]
  assign finder_1_io_data_5 = addrVec_5; // @[elements.scala 182:27]
  assign finder_1_io_data_6 = addrVec_6; // @[elements.scala 182:27]
  assign finder_1_io_data_7 = addrVec_7; // @[elements.scala 182:27]
  assign finder_1_io_data_8 = addrVec_8; // @[elements.scala 182:27]
  assign finder_1_io_data_9 = addrVec_9; // @[elements.scala 182:27]
  assign finder_1_io_data_10 = addrVec_10; // @[elements.scala 182:27]
  assign finder_1_io_data_11 = addrVec_11; // @[elements.scala 182:27]
  assign finder_1_io_data_12 = addrVec_12; // @[elements.scala 182:27]
  assign finder_1_io_data_13 = addrVec_13; // @[elements.scala 182:27]
  assign finder_1_io_data_14 = addrVec_14; // @[elements.scala 182:27]
  assign finder_1_io_data_15 = addrVec_15; // @[elements.scala 182:27]
  assign finder_1_io_valid_0 = valid_0; // @[elements.scala 184:28]
  assign finder_1_io_valid_1 = valid_1; // @[elements.scala 184:28]
  assign finder_1_io_valid_2 = valid_2; // @[elements.scala 184:28]
  assign finder_1_io_valid_3 = valid_3; // @[elements.scala 184:28]
  assign finder_1_io_valid_4 = valid_4; // @[elements.scala 184:28]
  assign finder_1_io_valid_5 = valid_5; // @[elements.scala 184:28]
  assign finder_1_io_valid_6 = valid_6; // @[elements.scala 184:28]
  assign finder_1_io_valid_7 = valid_7; // @[elements.scala 184:28]
  assign finder_1_io_valid_8 = valid_8; // @[elements.scala 184:28]
  assign finder_1_io_valid_9 = valid_9; // @[elements.scala 184:28]
  assign finder_1_io_valid_10 = valid_10; // @[elements.scala 184:28]
  assign finder_1_io_valid_11 = valid_11; // @[elements.scala 184:28]
  assign finder_1_io_valid_12 = valid_12; // @[elements.scala 184:28]
  assign finder_1_io_valid_13 = valid_13; // @[elements.scala 184:28]
  assign finder_1_io_valid_14 = valid_14; // @[elements.scala 184:28]
  assign finder_1_io_valid_15 = valid_15; // @[elements.scala 184:28]
  assign finder_2_io_key = io_unLock_2_in_bits_addr; // @[elements.scala 183:26]
  assign finder_2_io_data_0 = addrVec_0; // @[elements.scala 182:27]
  assign finder_2_io_data_1 = addrVec_1; // @[elements.scala 182:27]
  assign finder_2_io_data_2 = addrVec_2; // @[elements.scala 182:27]
  assign finder_2_io_data_3 = addrVec_3; // @[elements.scala 182:27]
  assign finder_2_io_data_4 = addrVec_4; // @[elements.scala 182:27]
  assign finder_2_io_data_5 = addrVec_5; // @[elements.scala 182:27]
  assign finder_2_io_data_6 = addrVec_6; // @[elements.scala 182:27]
  assign finder_2_io_data_7 = addrVec_7; // @[elements.scala 182:27]
  assign finder_2_io_data_8 = addrVec_8; // @[elements.scala 182:27]
  assign finder_2_io_data_9 = addrVec_9; // @[elements.scala 182:27]
  assign finder_2_io_data_10 = addrVec_10; // @[elements.scala 182:27]
  assign finder_2_io_data_11 = addrVec_11; // @[elements.scala 182:27]
  assign finder_2_io_data_12 = addrVec_12; // @[elements.scala 182:27]
  assign finder_2_io_data_13 = addrVec_13; // @[elements.scala 182:27]
  assign finder_2_io_data_14 = addrVec_14; // @[elements.scala 182:27]
  assign finder_2_io_data_15 = addrVec_15; // @[elements.scala 182:27]
  assign finder_2_io_valid_0 = valid_0; // @[elements.scala 184:28]
  assign finder_2_io_valid_1 = valid_1; // @[elements.scala 184:28]
  assign finder_2_io_valid_2 = valid_2; // @[elements.scala 184:28]
  assign finder_2_io_valid_3 = valid_3; // @[elements.scala 184:28]
  assign finder_2_io_valid_4 = valid_4; // @[elements.scala 184:28]
  assign finder_2_io_valid_5 = valid_5; // @[elements.scala 184:28]
  assign finder_2_io_valid_6 = valid_6; // @[elements.scala 184:28]
  assign finder_2_io_valid_7 = valid_7; // @[elements.scala 184:28]
  assign finder_2_io_valid_8 = valid_8; // @[elements.scala 184:28]
  assign finder_2_io_valid_9 = valid_9; // @[elements.scala 184:28]
  assign finder_2_io_valid_10 = valid_10; // @[elements.scala 184:28]
  assign finder_2_io_valid_11 = valid_11; // @[elements.scala 184:28]
  assign finder_2_io_valid_12 = valid_12; // @[elements.scala 184:28]
  assign finder_2_io_valid_13 = valid_13; // @[elements.scala 184:28]
  assign finder_2_io_valid_14 = valid_14; // @[elements.scala 184:28]
  assign finder_2_io_valid_15 = valid_15; // @[elements.scala 184:28]
  assign finder_3_io_key = io_unLock_3_in_bits_addr; // @[elements.scala 183:26]
  assign finder_3_io_data_0 = addrVec_0; // @[elements.scala 182:27]
  assign finder_3_io_data_1 = addrVec_1; // @[elements.scala 182:27]
  assign finder_3_io_data_2 = addrVec_2; // @[elements.scala 182:27]
  assign finder_3_io_data_3 = addrVec_3; // @[elements.scala 182:27]
  assign finder_3_io_data_4 = addrVec_4; // @[elements.scala 182:27]
  assign finder_3_io_data_5 = addrVec_5; // @[elements.scala 182:27]
  assign finder_3_io_data_6 = addrVec_6; // @[elements.scala 182:27]
  assign finder_3_io_data_7 = addrVec_7; // @[elements.scala 182:27]
  assign finder_3_io_data_8 = addrVec_8; // @[elements.scala 182:27]
  assign finder_3_io_data_9 = addrVec_9; // @[elements.scala 182:27]
  assign finder_3_io_data_10 = addrVec_10; // @[elements.scala 182:27]
  assign finder_3_io_data_11 = addrVec_11; // @[elements.scala 182:27]
  assign finder_3_io_data_12 = addrVec_12; // @[elements.scala 182:27]
  assign finder_3_io_data_13 = addrVec_13; // @[elements.scala 182:27]
  assign finder_3_io_data_14 = addrVec_14; // @[elements.scala 182:27]
  assign finder_3_io_data_15 = addrVec_15; // @[elements.scala 182:27]
  assign finder_3_io_valid_0 = valid_0; // @[elements.scala 184:28]
  assign finder_3_io_valid_1 = valid_1; // @[elements.scala 184:28]
  assign finder_3_io_valid_2 = valid_2; // @[elements.scala 184:28]
  assign finder_3_io_valid_3 = valid_3; // @[elements.scala 184:28]
  assign finder_3_io_valid_4 = valid_4; // @[elements.scala 184:28]
  assign finder_3_io_valid_5 = valid_5; // @[elements.scala 184:28]
  assign finder_3_io_valid_6 = valid_6; // @[elements.scala 184:28]
  assign finder_3_io_valid_7 = valid_7; // @[elements.scala 184:28]
  assign finder_3_io_valid_8 = valid_8; // @[elements.scala 184:28]
  assign finder_3_io_valid_9 = valid_9; // @[elements.scala 184:28]
  assign finder_3_io_valid_10 = valid_10; // @[elements.scala 184:28]
  assign finder_3_io_valid_11 = valid_11; // @[elements.scala 184:28]
  assign finder_3_io_valid_12 = valid_12; // @[elements.scala 184:28]
  assign finder_3_io_valid_13 = valid_13; // @[elements.scala 184:28]
  assign finder_3_io_valid_14 = valid_14; // @[elements.scala 184:28]
  assign finder_3_io_valid_15 = valid_15; // @[elements.scala 184:28]
  assign finder_4_io_key = io_unLock_4_in_bits_addr; // @[elements.scala 183:26]
  assign finder_4_io_data_0 = addrVec_0; // @[elements.scala 182:27]
  assign finder_4_io_data_1 = addrVec_1; // @[elements.scala 182:27]
  assign finder_4_io_data_2 = addrVec_2; // @[elements.scala 182:27]
  assign finder_4_io_data_3 = addrVec_3; // @[elements.scala 182:27]
  assign finder_4_io_data_4 = addrVec_4; // @[elements.scala 182:27]
  assign finder_4_io_data_5 = addrVec_5; // @[elements.scala 182:27]
  assign finder_4_io_data_6 = addrVec_6; // @[elements.scala 182:27]
  assign finder_4_io_data_7 = addrVec_7; // @[elements.scala 182:27]
  assign finder_4_io_data_8 = addrVec_8; // @[elements.scala 182:27]
  assign finder_4_io_data_9 = addrVec_9; // @[elements.scala 182:27]
  assign finder_4_io_data_10 = addrVec_10; // @[elements.scala 182:27]
  assign finder_4_io_data_11 = addrVec_11; // @[elements.scala 182:27]
  assign finder_4_io_data_12 = addrVec_12; // @[elements.scala 182:27]
  assign finder_4_io_data_13 = addrVec_13; // @[elements.scala 182:27]
  assign finder_4_io_data_14 = addrVec_14; // @[elements.scala 182:27]
  assign finder_4_io_data_15 = addrVec_15; // @[elements.scala 182:27]
  assign finder_4_io_valid_0 = valid_0; // @[elements.scala 184:28]
  assign finder_4_io_valid_1 = valid_1; // @[elements.scala 184:28]
  assign finder_4_io_valid_2 = valid_2; // @[elements.scala 184:28]
  assign finder_4_io_valid_3 = valid_3; // @[elements.scala 184:28]
  assign finder_4_io_valid_4 = valid_4; // @[elements.scala 184:28]
  assign finder_4_io_valid_5 = valid_5; // @[elements.scala 184:28]
  assign finder_4_io_valid_6 = valid_6; // @[elements.scala 184:28]
  assign finder_4_io_valid_7 = valid_7; // @[elements.scala 184:28]
  assign finder_4_io_valid_8 = valid_8; // @[elements.scala 184:28]
  assign finder_4_io_valid_9 = valid_9; // @[elements.scala 184:28]
  assign finder_4_io_valid_10 = valid_10; // @[elements.scala 184:28]
  assign finder_4_io_valid_11 = valid_11; // @[elements.scala 184:28]
  assign finder_4_io_valid_12 = valid_12; // @[elements.scala 184:28]
  assign finder_4_io_valid_13 = valid_13; // @[elements.scala 184:28]
  assign finder_4_io_valid_14 = valid_14; // @[elements.scala 184:28]
  assign finder_4_io_valid_15 = valid_15; // @[elements.scala 184:28]
  assign finder_5_io_key = io_unLock_5_in_bits_addr; // @[elements.scala 183:26]
  assign finder_5_io_data_0 = addrVec_0; // @[elements.scala 182:27]
  assign finder_5_io_data_1 = addrVec_1; // @[elements.scala 182:27]
  assign finder_5_io_data_2 = addrVec_2; // @[elements.scala 182:27]
  assign finder_5_io_data_3 = addrVec_3; // @[elements.scala 182:27]
  assign finder_5_io_data_4 = addrVec_4; // @[elements.scala 182:27]
  assign finder_5_io_data_5 = addrVec_5; // @[elements.scala 182:27]
  assign finder_5_io_data_6 = addrVec_6; // @[elements.scala 182:27]
  assign finder_5_io_data_7 = addrVec_7; // @[elements.scala 182:27]
  assign finder_5_io_data_8 = addrVec_8; // @[elements.scala 182:27]
  assign finder_5_io_data_9 = addrVec_9; // @[elements.scala 182:27]
  assign finder_5_io_data_10 = addrVec_10; // @[elements.scala 182:27]
  assign finder_5_io_data_11 = addrVec_11; // @[elements.scala 182:27]
  assign finder_5_io_data_12 = addrVec_12; // @[elements.scala 182:27]
  assign finder_5_io_data_13 = addrVec_13; // @[elements.scala 182:27]
  assign finder_5_io_data_14 = addrVec_14; // @[elements.scala 182:27]
  assign finder_5_io_data_15 = addrVec_15; // @[elements.scala 182:27]
  assign finder_5_io_valid_0 = valid_0; // @[elements.scala 184:28]
  assign finder_5_io_valid_1 = valid_1; // @[elements.scala 184:28]
  assign finder_5_io_valid_2 = valid_2; // @[elements.scala 184:28]
  assign finder_5_io_valid_3 = valid_3; // @[elements.scala 184:28]
  assign finder_5_io_valid_4 = valid_4; // @[elements.scala 184:28]
  assign finder_5_io_valid_5 = valid_5; // @[elements.scala 184:28]
  assign finder_5_io_valid_6 = valid_6; // @[elements.scala 184:28]
  assign finder_5_io_valid_7 = valid_7; // @[elements.scala 184:28]
  assign finder_5_io_valid_8 = valid_8; // @[elements.scala 184:28]
  assign finder_5_io_valid_9 = valid_9; // @[elements.scala 184:28]
  assign finder_5_io_valid_10 = valid_10; // @[elements.scala 184:28]
  assign finder_5_io_valid_11 = valid_11; // @[elements.scala 184:28]
  assign finder_5_io_valid_12 = valid_12; // @[elements.scala 184:28]
  assign finder_5_io_valid_13 = valid_13; // @[elements.scala 184:28]
  assign finder_5_io_valid_14 = valid_14; // @[elements.scala 184:28]
  assign finder_5_io_valid_15 = valid_15; // @[elements.scala 184:28]
  assign finder_6_io_key = io_unLock_6_in_bits_addr; // @[elements.scala 183:26]
  assign finder_6_io_data_0 = addrVec_0; // @[elements.scala 182:27]
  assign finder_6_io_data_1 = addrVec_1; // @[elements.scala 182:27]
  assign finder_6_io_data_2 = addrVec_2; // @[elements.scala 182:27]
  assign finder_6_io_data_3 = addrVec_3; // @[elements.scala 182:27]
  assign finder_6_io_data_4 = addrVec_4; // @[elements.scala 182:27]
  assign finder_6_io_data_5 = addrVec_5; // @[elements.scala 182:27]
  assign finder_6_io_data_6 = addrVec_6; // @[elements.scala 182:27]
  assign finder_6_io_data_7 = addrVec_7; // @[elements.scala 182:27]
  assign finder_6_io_data_8 = addrVec_8; // @[elements.scala 182:27]
  assign finder_6_io_data_9 = addrVec_9; // @[elements.scala 182:27]
  assign finder_6_io_data_10 = addrVec_10; // @[elements.scala 182:27]
  assign finder_6_io_data_11 = addrVec_11; // @[elements.scala 182:27]
  assign finder_6_io_data_12 = addrVec_12; // @[elements.scala 182:27]
  assign finder_6_io_data_13 = addrVec_13; // @[elements.scala 182:27]
  assign finder_6_io_data_14 = addrVec_14; // @[elements.scala 182:27]
  assign finder_6_io_data_15 = addrVec_15; // @[elements.scala 182:27]
  assign finder_6_io_valid_0 = valid_0; // @[elements.scala 184:28]
  assign finder_6_io_valid_1 = valid_1; // @[elements.scala 184:28]
  assign finder_6_io_valid_2 = valid_2; // @[elements.scala 184:28]
  assign finder_6_io_valid_3 = valid_3; // @[elements.scala 184:28]
  assign finder_6_io_valid_4 = valid_4; // @[elements.scala 184:28]
  assign finder_6_io_valid_5 = valid_5; // @[elements.scala 184:28]
  assign finder_6_io_valid_6 = valid_6; // @[elements.scala 184:28]
  assign finder_6_io_valid_7 = valid_7; // @[elements.scala 184:28]
  assign finder_6_io_valid_8 = valid_8; // @[elements.scala 184:28]
  assign finder_6_io_valid_9 = valid_9; // @[elements.scala 184:28]
  assign finder_6_io_valid_10 = valid_10; // @[elements.scala 184:28]
  assign finder_6_io_valid_11 = valid_11; // @[elements.scala 184:28]
  assign finder_6_io_valid_12 = valid_12; // @[elements.scala 184:28]
  assign finder_6_io_valid_13 = valid_13; // @[elements.scala 184:28]
  assign finder_6_io_valid_14 = valid_14; // @[elements.scala 184:28]
  assign finder_6_io_valid_15 = valid_15; // @[elements.scala 184:28]
  assign finder_7_io_key = io_unLock_7_in_bits_addr; // @[elements.scala 183:26]
  assign finder_7_io_data_0 = addrVec_0; // @[elements.scala 182:27]
  assign finder_7_io_data_1 = addrVec_1; // @[elements.scala 182:27]
  assign finder_7_io_data_2 = addrVec_2; // @[elements.scala 182:27]
  assign finder_7_io_data_3 = addrVec_3; // @[elements.scala 182:27]
  assign finder_7_io_data_4 = addrVec_4; // @[elements.scala 182:27]
  assign finder_7_io_data_5 = addrVec_5; // @[elements.scala 182:27]
  assign finder_7_io_data_6 = addrVec_6; // @[elements.scala 182:27]
  assign finder_7_io_data_7 = addrVec_7; // @[elements.scala 182:27]
  assign finder_7_io_data_8 = addrVec_8; // @[elements.scala 182:27]
  assign finder_7_io_data_9 = addrVec_9; // @[elements.scala 182:27]
  assign finder_7_io_data_10 = addrVec_10; // @[elements.scala 182:27]
  assign finder_7_io_data_11 = addrVec_11; // @[elements.scala 182:27]
  assign finder_7_io_data_12 = addrVec_12; // @[elements.scala 182:27]
  assign finder_7_io_data_13 = addrVec_13; // @[elements.scala 182:27]
  assign finder_7_io_data_14 = addrVec_14; // @[elements.scala 182:27]
  assign finder_7_io_data_15 = addrVec_15; // @[elements.scala 182:27]
  assign finder_7_io_valid_0 = valid_0; // @[elements.scala 184:28]
  assign finder_7_io_valid_1 = valid_1; // @[elements.scala 184:28]
  assign finder_7_io_valid_2 = valid_2; // @[elements.scala 184:28]
  assign finder_7_io_valid_3 = valid_3; // @[elements.scala 184:28]
  assign finder_7_io_valid_4 = valid_4; // @[elements.scala 184:28]
  assign finder_7_io_valid_5 = valid_5; // @[elements.scala 184:28]
  assign finder_7_io_valid_6 = valid_6; // @[elements.scala 184:28]
  assign finder_7_io_valid_7 = valid_7; // @[elements.scala 184:28]
  assign finder_7_io_valid_8 = valid_8; // @[elements.scala 184:28]
  assign finder_7_io_valid_9 = valid_9; // @[elements.scala 184:28]
  assign finder_7_io_valid_10 = valid_10; // @[elements.scala 184:28]
  assign finder_7_io_valid_11 = valid_11; // @[elements.scala 184:28]
  assign finder_7_io_valid_12 = valid_12; // @[elements.scala 184:28]
  assign finder_7_io_valid_13 = valid_13; // @[elements.scala 184:28]
  assign finder_7_io_valid_14 = valid_14; // @[elements.scala 184:28]
  assign finder_7_io_valid_15 = valid_15; // @[elements.scala 184:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addrVec_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  addrVec_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  addrVec_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  addrVec_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  addrVec_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  addrVec_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  addrVec_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  addrVec_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  addrVec_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  addrVec_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  addrVec_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  addrVec_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  addrVec_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  addrVec_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  addrVec_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  addrVec_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  valid_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_4 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_5 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_6 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_7 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_8 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_9 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_10 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_11 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_12 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_13 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_14 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_15 = _RAND_31[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addrVec_0 <= 32'h0;
    end else if (write) begin
      if (4'h0 == idxLocking[3:0]) begin
        addrVec_0 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_1 <= 32'h0;
    end else if (write) begin
      if (4'h1 == idxLocking[3:0]) begin
        addrVec_1 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_2 <= 32'h0;
    end else if (write) begin
      if (4'h2 == idxLocking[3:0]) begin
        addrVec_2 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_3 <= 32'h0;
    end else if (write) begin
      if (4'h3 == idxLocking[3:0]) begin
        addrVec_3 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_4 <= 32'h0;
    end else if (write) begin
      if (4'h4 == idxLocking[3:0]) begin
        addrVec_4 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_5 <= 32'h0;
    end else if (write) begin
      if (4'h5 == idxLocking[3:0]) begin
        addrVec_5 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_6 <= 32'h0;
    end else if (write) begin
      if (4'h6 == idxLocking[3:0]) begin
        addrVec_6 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_7 <= 32'h0;
    end else if (write) begin
      if (4'h7 == idxLocking[3:0]) begin
        addrVec_7 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_8 <= 32'h0;
    end else if (write) begin
      if (4'h8 == idxLocking[3:0]) begin
        addrVec_8 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_9 <= 32'h0;
    end else if (write) begin
      if (4'h9 == idxLocking[3:0]) begin
        addrVec_9 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_10 <= 32'h0;
    end else if (write) begin
      if (4'ha == idxLocking[3:0]) begin
        addrVec_10 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_11 <= 32'h0;
    end else if (write) begin
      if (4'hb == idxLocking[3:0]) begin
        addrVec_11 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_12 <= 32'h0;
    end else if (write) begin
      if (4'hc == idxLocking[3:0]) begin
        addrVec_12 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_13 <= 32'h0;
    end else if (write) begin
      if (4'hd == idxLocking[3:0]) begin
        addrVec_13 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_14 <= 32'h0;
    end else if (write) begin
      if (4'he == idxLocking[3:0]) begin
        addrVec_14 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      addrVec_15 <= 32'h0;
    end else if (write) begin
      if (4'hf == idxLocking[3:0]) begin
        addrVec_15 <= io_lock_in_bits_addr;
      end
    end
    if (reset) begin
      valid_0 <= 1'h0;
    end else if (write) begin
      valid_0 <= _GEN_305;
    end else if (_T_125) begin
      if (4'h0 == idxUnlock_7[3:0]) begin
        valid_0 <= 1'h0;
      end else if (_T_123) begin
        if (4'h0 == idxUnlock_6[3:0]) begin
          valid_0 <= 1'h0;
        end else if (_T_121) begin
          if (4'h0 == idxUnlock_5[3:0]) begin
            valid_0 <= 1'h0;
          end else if (_T_119) begin
            if (4'h0 == idxUnlock_4[3:0]) begin
              valid_0 <= 1'h0;
            end else if (_T_117) begin
              if (4'h0 == idxUnlock_3[3:0]) begin
                valid_0 <= 1'h0;
              end else if (_T_115) begin
                if (4'h0 == idxUnlock_2[3:0]) begin
                  valid_0 <= 1'h0;
                end else if (_T_113) begin
                  if (4'h0 == idxUnlock_1[3:0]) begin
                    valid_0 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'h0 == idxUnlock_0[3:0]) begin
                      valid_0 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h0 == idxUnlock_0[3:0]) begin
                    valid_0 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'h0 == idxUnlock_1[3:0]) begin
                  valid_0 <= 1'h0;
                end else if (_T_111) begin
                  if (4'h0 == idxUnlock_0[3:0]) begin
                    valid_0 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'h0 == idxUnlock_0[3:0]) begin
                  valid_0 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'h0 == idxUnlock_2[3:0]) begin
                valid_0 <= 1'h0;
              end else if (_T_113) begin
                if (4'h0 == idxUnlock_1[3:0]) begin
                  valid_0 <= 1'h0;
                end else begin
                  valid_0 <= _GEN_16;
                end
              end else begin
                valid_0 <= _GEN_16;
              end
            end else if (_T_113) begin
              if (4'h0 == idxUnlock_1[3:0]) begin
                valid_0 <= 1'h0;
              end else begin
                valid_0 <= _GEN_16;
              end
            end else begin
              valid_0 <= _GEN_16;
            end
          end else if (_T_117) begin
            if (4'h0 == idxUnlock_3[3:0]) begin
              valid_0 <= 1'h0;
            end else if (_T_115) begin
              if (4'h0 == idxUnlock_2[3:0]) begin
                valid_0 <= 1'h0;
              end else begin
                valid_0 <= _GEN_48;
              end
            end else begin
              valid_0 <= _GEN_48;
            end
          end else if (_T_115) begin
            if (4'h0 == idxUnlock_2[3:0]) begin
              valid_0 <= 1'h0;
            end else begin
              valid_0 <= _GEN_48;
            end
          end else begin
            valid_0 <= _GEN_48;
          end
        end else if (_T_119) begin
          if (4'h0 == idxUnlock_4[3:0]) begin
            valid_0 <= 1'h0;
          end else if (_T_117) begin
            if (4'h0 == idxUnlock_3[3:0]) begin
              valid_0 <= 1'h0;
            end else begin
              valid_0 <= _GEN_80;
            end
          end else begin
            valid_0 <= _GEN_80;
          end
        end else if (_T_117) begin
          if (4'h0 == idxUnlock_3[3:0]) begin
            valid_0 <= 1'h0;
          end else begin
            valid_0 <= _GEN_80;
          end
        end else begin
          valid_0 <= _GEN_80;
        end
      end else if (_T_121) begin
        if (4'h0 == idxUnlock_5[3:0]) begin
          valid_0 <= 1'h0;
        end else if (_T_119) begin
          if (4'h0 == idxUnlock_4[3:0]) begin
            valid_0 <= 1'h0;
          end else begin
            valid_0 <= _GEN_112;
          end
        end else begin
          valid_0 <= _GEN_112;
        end
      end else if (_T_119) begin
        if (4'h0 == idxUnlock_4[3:0]) begin
          valid_0 <= 1'h0;
        end else begin
          valid_0 <= _GEN_112;
        end
      end else begin
        valid_0 <= _GEN_112;
      end
    end else if (_T_123) begin
      if (4'h0 == idxUnlock_6[3:0]) begin
        valid_0 <= 1'h0;
      end else if (_T_121) begin
        if (4'h0 == idxUnlock_5[3:0]) begin
          valid_0 <= 1'h0;
        end else begin
          valid_0 <= _GEN_144;
        end
      end else begin
        valid_0 <= _GEN_144;
      end
    end else if (_T_121) begin
      if (4'h0 == idxUnlock_5[3:0]) begin
        valid_0 <= 1'h0;
      end else begin
        valid_0 <= _GEN_144;
      end
    end else begin
      valid_0 <= _GEN_144;
    end
    if (reset) begin
      valid_1 <= 1'h0;
    end else if (write) begin
      valid_1 <= _GEN_306;
    end else if (_T_125) begin
      if (4'h1 == idxUnlock_7[3:0]) begin
        valid_1 <= 1'h0;
      end else if (_T_123) begin
        if (4'h1 == idxUnlock_6[3:0]) begin
          valid_1 <= 1'h0;
        end else if (_T_121) begin
          if (4'h1 == idxUnlock_5[3:0]) begin
            valid_1 <= 1'h0;
          end else if (_T_119) begin
            if (4'h1 == idxUnlock_4[3:0]) begin
              valid_1 <= 1'h0;
            end else if (_T_117) begin
              if (4'h1 == idxUnlock_3[3:0]) begin
                valid_1 <= 1'h0;
              end else if (_T_115) begin
                if (4'h1 == idxUnlock_2[3:0]) begin
                  valid_1 <= 1'h0;
                end else if (_T_113) begin
                  if (4'h1 == idxUnlock_1[3:0]) begin
                    valid_1 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'h1 == idxUnlock_0[3:0]) begin
                      valid_1 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h1 == idxUnlock_0[3:0]) begin
                    valid_1 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'h1 == idxUnlock_1[3:0]) begin
                  valid_1 <= 1'h0;
                end else if (_T_111) begin
                  if (4'h1 == idxUnlock_0[3:0]) begin
                    valid_1 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'h1 == idxUnlock_0[3:0]) begin
                  valid_1 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'h1 == idxUnlock_2[3:0]) begin
                valid_1 <= 1'h0;
              end else if (_T_113) begin
                if (4'h1 == idxUnlock_1[3:0]) begin
                  valid_1 <= 1'h0;
                end else begin
                  valid_1 <= _GEN_17;
                end
              end else begin
                valid_1 <= _GEN_17;
              end
            end else if (_T_113) begin
              if (4'h1 == idxUnlock_1[3:0]) begin
                valid_1 <= 1'h0;
              end else begin
                valid_1 <= _GEN_17;
              end
            end else begin
              valid_1 <= _GEN_17;
            end
          end else if (_T_117) begin
            if (4'h1 == idxUnlock_3[3:0]) begin
              valid_1 <= 1'h0;
            end else if (_T_115) begin
              if (4'h1 == idxUnlock_2[3:0]) begin
                valid_1 <= 1'h0;
              end else begin
                valid_1 <= _GEN_49;
              end
            end else begin
              valid_1 <= _GEN_49;
            end
          end else if (_T_115) begin
            if (4'h1 == idxUnlock_2[3:0]) begin
              valid_1 <= 1'h0;
            end else begin
              valid_1 <= _GEN_49;
            end
          end else begin
            valid_1 <= _GEN_49;
          end
        end else if (_T_119) begin
          if (4'h1 == idxUnlock_4[3:0]) begin
            valid_1 <= 1'h0;
          end else if (_T_117) begin
            if (4'h1 == idxUnlock_3[3:0]) begin
              valid_1 <= 1'h0;
            end else begin
              valid_1 <= _GEN_81;
            end
          end else begin
            valid_1 <= _GEN_81;
          end
        end else if (_T_117) begin
          if (4'h1 == idxUnlock_3[3:0]) begin
            valid_1 <= 1'h0;
          end else begin
            valid_1 <= _GEN_81;
          end
        end else begin
          valid_1 <= _GEN_81;
        end
      end else if (_T_121) begin
        if (4'h1 == idxUnlock_5[3:0]) begin
          valid_1 <= 1'h0;
        end else if (_T_119) begin
          if (4'h1 == idxUnlock_4[3:0]) begin
            valid_1 <= 1'h0;
          end else begin
            valid_1 <= _GEN_113;
          end
        end else begin
          valid_1 <= _GEN_113;
        end
      end else if (_T_119) begin
        if (4'h1 == idxUnlock_4[3:0]) begin
          valid_1 <= 1'h0;
        end else begin
          valid_1 <= _GEN_113;
        end
      end else begin
        valid_1 <= _GEN_113;
      end
    end else if (_T_123) begin
      if (4'h1 == idxUnlock_6[3:0]) begin
        valid_1 <= 1'h0;
      end else if (_T_121) begin
        if (4'h1 == idxUnlock_5[3:0]) begin
          valid_1 <= 1'h0;
        end else begin
          valid_1 <= _GEN_145;
        end
      end else begin
        valid_1 <= _GEN_145;
      end
    end else if (_T_121) begin
      if (4'h1 == idxUnlock_5[3:0]) begin
        valid_1 <= 1'h0;
      end else begin
        valid_1 <= _GEN_145;
      end
    end else begin
      valid_1 <= _GEN_145;
    end
    if (reset) begin
      valid_2 <= 1'h0;
    end else if (write) begin
      valid_2 <= _GEN_307;
    end else if (_T_125) begin
      if (4'h2 == idxUnlock_7[3:0]) begin
        valid_2 <= 1'h0;
      end else if (_T_123) begin
        if (4'h2 == idxUnlock_6[3:0]) begin
          valid_2 <= 1'h0;
        end else if (_T_121) begin
          if (4'h2 == idxUnlock_5[3:0]) begin
            valid_2 <= 1'h0;
          end else if (_T_119) begin
            if (4'h2 == idxUnlock_4[3:0]) begin
              valid_2 <= 1'h0;
            end else if (_T_117) begin
              if (4'h2 == idxUnlock_3[3:0]) begin
                valid_2 <= 1'h0;
              end else if (_T_115) begin
                if (4'h2 == idxUnlock_2[3:0]) begin
                  valid_2 <= 1'h0;
                end else if (_T_113) begin
                  if (4'h2 == idxUnlock_1[3:0]) begin
                    valid_2 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'h2 == idxUnlock_0[3:0]) begin
                      valid_2 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h2 == idxUnlock_0[3:0]) begin
                    valid_2 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'h2 == idxUnlock_1[3:0]) begin
                  valid_2 <= 1'h0;
                end else if (_T_111) begin
                  if (4'h2 == idxUnlock_0[3:0]) begin
                    valid_2 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'h2 == idxUnlock_0[3:0]) begin
                  valid_2 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'h2 == idxUnlock_2[3:0]) begin
                valid_2 <= 1'h0;
              end else if (_T_113) begin
                if (4'h2 == idxUnlock_1[3:0]) begin
                  valid_2 <= 1'h0;
                end else begin
                  valid_2 <= _GEN_18;
                end
              end else begin
                valid_2 <= _GEN_18;
              end
            end else if (_T_113) begin
              if (4'h2 == idxUnlock_1[3:0]) begin
                valid_2 <= 1'h0;
              end else begin
                valid_2 <= _GEN_18;
              end
            end else begin
              valid_2 <= _GEN_18;
            end
          end else if (_T_117) begin
            if (4'h2 == idxUnlock_3[3:0]) begin
              valid_2 <= 1'h0;
            end else if (_T_115) begin
              if (4'h2 == idxUnlock_2[3:0]) begin
                valid_2 <= 1'h0;
              end else begin
                valid_2 <= _GEN_50;
              end
            end else begin
              valid_2 <= _GEN_50;
            end
          end else if (_T_115) begin
            if (4'h2 == idxUnlock_2[3:0]) begin
              valid_2 <= 1'h0;
            end else begin
              valid_2 <= _GEN_50;
            end
          end else begin
            valid_2 <= _GEN_50;
          end
        end else if (_T_119) begin
          if (4'h2 == idxUnlock_4[3:0]) begin
            valid_2 <= 1'h0;
          end else if (_T_117) begin
            if (4'h2 == idxUnlock_3[3:0]) begin
              valid_2 <= 1'h0;
            end else begin
              valid_2 <= _GEN_82;
            end
          end else begin
            valid_2 <= _GEN_82;
          end
        end else if (_T_117) begin
          if (4'h2 == idxUnlock_3[3:0]) begin
            valid_2 <= 1'h0;
          end else begin
            valid_2 <= _GEN_82;
          end
        end else begin
          valid_2 <= _GEN_82;
        end
      end else if (_T_121) begin
        if (4'h2 == idxUnlock_5[3:0]) begin
          valid_2 <= 1'h0;
        end else if (_T_119) begin
          if (4'h2 == idxUnlock_4[3:0]) begin
            valid_2 <= 1'h0;
          end else begin
            valid_2 <= _GEN_114;
          end
        end else begin
          valid_2 <= _GEN_114;
        end
      end else if (_T_119) begin
        if (4'h2 == idxUnlock_4[3:0]) begin
          valid_2 <= 1'h0;
        end else begin
          valid_2 <= _GEN_114;
        end
      end else begin
        valid_2 <= _GEN_114;
      end
    end else if (_T_123) begin
      if (4'h2 == idxUnlock_6[3:0]) begin
        valid_2 <= 1'h0;
      end else if (_T_121) begin
        if (4'h2 == idxUnlock_5[3:0]) begin
          valid_2 <= 1'h0;
        end else begin
          valid_2 <= _GEN_146;
        end
      end else begin
        valid_2 <= _GEN_146;
      end
    end else if (_T_121) begin
      if (4'h2 == idxUnlock_5[3:0]) begin
        valid_2 <= 1'h0;
      end else begin
        valid_2 <= _GEN_146;
      end
    end else begin
      valid_2 <= _GEN_146;
    end
    if (reset) begin
      valid_3 <= 1'h0;
    end else if (write) begin
      valid_3 <= _GEN_308;
    end else if (_T_125) begin
      if (4'h3 == idxUnlock_7[3:0]) begin
        valid_3 <= 1'h0;
      end else if (_T_123) begin
        if (4'h3 == idxUnlock_6[3:0]) begin
          valid_3 <= 1'h0;
        end else if (_T_121) begin
          if (4'h3 == idxUnlock_5[3:0]) begin
            valid_3 <= 1'h0;
          end else if (_T_119) begin
            if (4'h3 == idxUnlock_4[3:0]) begin
              valid_3 <= 1'h0;
            end else if (_T_117) begin
              if (4'h3 == idxUnlock_3[3:0]) begin
                valid_3 <= 1'h0;
              end else if (_T_115) begin
                if (4'h3 == idxUnlock_2[3:0]) begin
                  valid_3 <= 1'h0;
                end else if (_T_113) begin
                  if (4'h3 == idxUnlock_1[3:0]) begin
                    valid_3 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'h3 == idxUnlock_0[3:0]) begin
                      valid_3 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h3 == idxUnlock_0[3:0]) begin
                    valid_3 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'h3 == idxUnlock_1[3:0]) begin
                  valid_3 <= 1'h0;
                end else if (_T_111) begin
                  if (4'h3 == idxUnlock_0[3:0]) begin
                    valid_3 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'h3 == idxUnlock_0[3:0]) begin
                  valid_3 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'h3 == idxUnlock_2[3:0]) begin
                valid_3 <= 1'h0;
              end else if (_T_113) begin
                if (4'h3 == idxUnlock_1[3:0]) begin
                  valid_3 <= 1'h0;
                end else begin
                  valid_3 <= _GEN_19;
                end
              end else begin
                valid_3 <= _GEN_19;
              end
            end else if (_T_113) begin
              if (4'h3 == idxUnlock_1[3:0]) begin
                valid_3 <= 1'h0;
              end else begin
                valid_3 <= _GEN_19;
              end
            end else begin
              valid_3 <= _GEN_19;
            end
          end else if (_T_117) begin
            if (4'h3 == idxUnlock_3[3:0]) begin
              valid_3 <= 1'h0;
            end else if (_T_115) begin
              if (4'h3 == idxUnlock_2[3:0]) begin
                valid_3 <= 1'h0;
              end else begin
                valid_3 <= _GEN_51;
              end
            end else begin
              valid_3 <= _GEN_51;
            end
          end else if (_T_115) begin
            if (4'h3 == idxUnlock_2[3:0]) begin
              valid_3 <= 1'h0;
            end else begin
              valid_3 <= _GEN_51;
            end
          end else begin
            valid_3 <= _GEN_51;
          end
        end else if (_T_119) begin
          if (4'h3 == idxUnlock_4[3:0]) begin
            valid_3 <= 1'h0;
          end else if (_T_117) begin
            if (4'h3 == idxUnlock_3[3:0]) begin
              valid_3 <= 1'h0;
            end else begin
              valid_3 <= _GEN_83;
            end
          end else begin
            valid_3 <= _GEN_83;
          end
        end else if (_T_117) begin
          if (4'h3 == idxUnlock_3[3:0]) begin
            valid_3 <= 1'h0;
          end else begin
            valid_3 <= _GEN_83;
          end
        end else begin
          valid_3 <= _GEN_83;
        end
      end else if (_T_121) begin
        if (4'h3 == idxUnlock_5[3:0]) begin
          valid_3 <= 1'h0;
        end else if (_T_119) begin
          if (4'h3 == idxUnlock_4[3:0]) begin
            valid_3 <= 1'h0;
          end else begin
            valid_3 <= _GEN_115;
          end
        end else begin
          valid_3 <= _GEN_115;
        end
      end else if (_T_119) begin
        if (4'h3 == idxUnlock_4[3:0]) begin
          valid_3 <= 1'h0;
        end else begin
          valid_3 <= _GEN_115;
        end
      end else begin
        valid_3 <= _GEN_115;
      end
    end else if (_T_123) begin
      if (4'h3 == idxUnlock_6[3:0]) begin
        valid_3 <= 1'h0;
      end else if (_T_121) begin
        if (4'h3 == idxUnlock_5[3:0]) begin
          valid_3 <= 1'h0;
        end else begin
          valid_3 <= _GEN_147;
        end
      end else begin
        valid_3 <= _GEN_147;
      end
    end else if (_T_121) begin
      if (4'h3 == idxUnlock_5[3:0]) begin
        valid_3 <= 1'h0;
      end else begin
        valid_3 <= _GEN_147;
      end
    end else begin
      valid_3 <= _GEN_147;
    end
    if (reset) begin
      valid_4 <= 1'h0;
    end else if (write) begin
      valid_4 <= _GEN_309;
    end else if (_T_125) begin
      if (4'h4 == idxUnlock_7[3:0]) begin
        valid_4 <= 1'h0;
      end else if (_T_123) begin
        if (4'h4 == idxUnlock_6[3:0]) begin
          valid_4 <= 1'h0;
        end else if (_T_121) begin
          if (4'h4 == idxUnlock_5[3:0]) begin
            valid_4 <= 1'h0;
          end else if (_T_119) begin
            if (4'h4 == idxUnlock_4[3:0]) begin
              valid_4 <= 1'h0;
            end else if (_T_117) begin
              if (4'h4 == idxUnlock_3[3:0]) begin
                valid_4 <= 1'h0;
              end else if (_T_115) begin
                if (4'h4 == idxUnlock_2[3:0]) begin
                  valid_4 <= 1'h0;
                end else if (_T_113) begin
                  if (4'h4 == idxUnlock_1[3:0]) begin
                    valid_4 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'h4 == idxUnlock_0[3:0]) begin
                      valid_4 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h4 == idxUnlock_0[3:0]) begin
                    valid_4 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'h4 == idxUnlock_1[3:0]) begin
                  valid_4 <= 1'h0;
                end else if (_T_111) begin
                  if (4'h4 == idxUnlock_0[3:0]) begin
                    valid_4 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'h4 == idxUnlock_0[3:0]) begin
                  valid_4 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'h4 == idxUnlock_2[3:0]) begin
                valid_4 <= 1'h0;
              end else if (_T_113) begin
                if (4'h4 == idxUnlock_1[3:0]) begin
                  valid_4 <= 1'h0;
                end else begin
                  valid_4 <= _GEN_20;
                end
              end else begin
                valid_4 <= _GEN_20;
              end
            end else if (_T_113) begin
              if (4'h4 == idxUnlock_1[3:0]) begin
                valid_4 <= 1'h0;
              end else begin
                valid_4 <= _GEN_20;
              end
            end else begin
              valid_4 <= _GEN_20;
            end
          end else if (_T_117) begin
            if (4'h4 == idxUnlock_3[3:0]) begin
              valid_4 <= 1'h0;
            end else if (_T_115) begin
              if (4'h4 == idxUnlock_2[3:0]) begin
                valid_4 <= 1'h0;
              end else begin
                valid_4 <= _GEN_52;
              end
            end else begin
              valid_4 <= _GEN_52;
            end
          end else if (_T_115) begin
            if (4'h4 == idxUnlock_2[3:0]) begin
              valid_4 <= 1'h0;
            end else begin
              valid_4 <= _GEN_52;
            end
          end else begin
            valid_4 <= _GEN_52;
          end
        end else if (_T_119) begin
          if (4'h4 == idxUnlock_4[3:0]) begin
            valid_4 <= 1'h0;
          end else if (_T_117) begin
            if (4'h4 == idxUnlock_3[3:0]) begin
              valid_4 <= 1'h0;
            end else begin
              valid_4 <= _GEN_84;
            end
          end else begin
            valid_4 <= _GEN_84;
          end
        end else if (_T_117) begin
          if (4'h4 == idxUnlock_3[3:0]) begin
            valid_4 <= 1'h0;
          end else begin
            valid_4 <= _GEN_84;
          end
        end else begin
          valid_4 <= _GEN_84;
        end
      end else if (_T_121) begin
        if (4'h4 == idxUnlock_5[3:0]) begin
          valid_4 <= 1'h0;
        end else if (_T_119) begin
          if (4'h4 == idxUnlock_4[3:0]) begin
            valid_4 <= 1'h0;
          end else begin
            valid_4 <= _GEN_116;
          end
        end else begin
          valid_4 <= _GEN_116;
        end
      end else if (_T_119) begin
        if (4'h4 == idxUnlock_4[3:0]) begin
          valid_4 <= 1'h0;
        end else begin
          valid_4 <= _GEN_116;
        end
      end else begin
        valid_4 <= _GEN_116;
      end
    end else if (_T_123) begin
      if (4'h4 == idxUnlock_6[3:0]) begin
        valid_4 <= 1'h0;
      end else if (_T_121) begin
        if (4'h4 == idxUnlock_5[3:0]) begin
          valid_4 <= 1'h0;
        end else begin
          valid_4 <= _GEN_148;
        end
      end else begin
        valid_4 <= _GEN_148;
      end
    end else if (_T_121) begin
      if (4'h4 == idxUnlock_5[3:0]) begin
        valid_4 <= 1'h0;
      end else begin
        valid_4 <= _GEN_148;
      end
    end else begin
      valid_4 <= _GEN_148;
    end
    if (reset) begin
      valid_5 <= 1'h0;
    end else if (write) begin
      valid_5 <= _GEN_310;
    end else if (_T_125) begin
      if (4'h5 == idxUnlock_7[3:0]) begin
        valid_5 <= 1'h0;
      end else if (_T_123) begin
        if (4'h5 == idxUnlock_6[3:0]) begin
          valid_5 <= 1'h0;
        end else if (_T_121) begin
          if (4'h5 == idxUnlock_5[3:0]) begin
            valid_5 <= 1'h0;
          end else if (_T_119) begin
            if (4'h5 == idxUnlock_4[3:0]) begin
              valid_5 <= 1'h0;
            end else if (_T_117) begin
              if (4'h5 == idxUnlock_3[3:0]) begin
                valid_5 <= 1'h0;
              end else if (_T_115) begin
                if (4'h5 == idxUnlock_2[3:0]) begin
                  valid_5 <= 1'h0;
                end else if (_T_113) begin
                  if (4'h5 == idxUnlock_1[3:0]) begin
                    valid_5 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'h5 == idxUnlock_0[3:0]) begin
                      valid_5 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h5 == idxUnlock_0[3:0]) begin
                    valid_5 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'h5 == idxUnlock_1[3:0]) begin
                  valid_5 <= 1'h0;
                end else if (_T_111) begin
                  if (4'h5 == idxUnlock_0[3:0]) begin
                    valid_5 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'h5 == idxUnlock_0[3:0]) begin
                  valid_5 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'h5 == idxUnlock_2[3:0]) begin
                valid_5 <= 1'h0;
              end else if (_T_113) begin
                if (4'h5 == idxUnlock_1[3:0]) begin
                  valid_5 <= 1'h0;
                end else begin
                  valid_5 <= _GEN_21;
                end
              end else begin
                valid_5 <= _GEN_21;
              end
            end else if (_T_113) begin
              if (4'h5 == idxUnlock_1[3:0]) begin
                valid_5 <= 1'h0;
              end else begin
                valid_5 <= _GEN_21;
              end
            end else begin
              valid_5 <= _GEN_21;
            end
          end else if (_T_117) begin
            if (4'h5 == idxUnlock_3[3:0]) begin
              valid_5 <= 1'h0;
            end else if (_T_115) begin
              if (4'h5 == idxUnlock_2[3:0]) begin
                valid_5 <= 1'h0;
              end else begin
                valid_5 <= _GEN_53;
              end
            end else begin
              valid_5 <= _GEN_53;
            end
          end else if (_T_115) begin
            if (4'h5 == idxUnlock_2[3:0]) begin
              valid_5 <= 1'h0;
            end else begin
              valid_5 <= _GEN_53;
            end
          end else begin
            valid_5 <= _GEN_53;
          end
        end else if (_T_119) begin
          if (4'h5 == idxUnlock_4[3:0]) begin
            valid_5 <= 1'h0;
          end else if (_T_117) begin
            if (4'h5 == idxUnlock_3[3:0]) begin
              valid_5 <= 1'h0;
            end else begin
              valid_5 <= _GEN_85;
            end
          end else begin
            valid_5 <= _GEN_85;
          end
        end else if (_T_117) begin
          if (4'h5 == idxUnlock_3[3:0]) begin
            valid_5 <= 1'h0;
          end else begin
            valid_5 <= _GEN_85;
          end
        end else begin
          valid_5 <= _GEN_85;
        end
      end else if (_T_121) begin
        if (4'h5 == idxUnlock_5[3:0]) begin
          valid_5 <= 1'h0;
        end else if (_T_119) begin
          if (4'h5 == idxUnlock_4[3:0]) begin
            valid_5 <= 1'h0;
          end else begin
            valid_5 <= _GEN_117;
          end
        end else begin
          valid_5 <= _GEN_117;
        end
      end else if (_T_119) begin
        if (4'h5 == idxUnlock_4[3:0]) begin
          valid_5 <= 1'h0;
        end else begin
          valid_5 <= _GEN_117;
        end
      end else begin
        valid_5 <= _GEN_117;
      end
    end else if (_T_123) begin
      if (4'h5 == idxUnlock_6[3:0]) begin
        valid_5 <= 1'h0;
      end else if (_T_121) begin
        if (4'h5 == idxUnlock_5[3:0]) begin
          valid_5 <= 1'h0;
        end else begin
          valid_5 <= _GEN_149;
        end
      end else begin
        valid_5 <= _GEN_149;
      end
    end else if (_T_121) begin
      if (4'h5 == idxUnlock_5[3:0]) begin
        valid_5 <= 1'h0;
      end else begin
        valid_5 <= _GEN_149;
      end
    end else begin
      valid_5 <= _GEN_149;
    end
    if (reset) begin
      valid_6 <= 1'h0;
    end else if (write) begin
      valid_6 <= _GEN_311;
    end else if (_T_125) begin
      if (4'h6 == idxUnlock_7[3:0]) begin
        valid_6 <= 1'h0;
      end else if (_T_123) begin
        if (4'h6 == idxUnlock_6[3:0]) begin
          valid_6 <= 1'h0;
        end else if (_T_121) begin
          if (4'h6 == idxUnlock_5[3:0]) begin
            valid_6 <= 1'h0;
          end else if (_T_119) begin
            if (4'h6 == idxUnlock_4[3:0]) begin
              valid_6 <= 1'h0;
            end else if (_T_117) begin
              if (4'h6 == idxUnlock_3[3:0]) begin
                valid_6 <= 1'h0;
              end else if (_T_115) begin
                if (4'h6 == idxUnlock_2[3:0]) begin
                  valid_6 <= 1'h0;
                end else if (_T_113) begin
                  if (4'h6 == idxUnlock_1[3:0]) begin
                    valid_6 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'h6 == idxUnlock_0[3:0]) begin
                      valid_6 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h6 == idxUnlock_0[3:0]) begin
                    valid_6 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'h6 == idxUnlock_1[3:0]) begin
                  valid_6 <= 1'h0;
                end else if (_T_111) begin
                  if (4'h6 == idxUnlock_0[3:0]) begin
                    valid_6 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'h6 == idxUnlock_0[3:0]) begin
                  valid_6 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'h6 == idxUnlock_2[3:0]) begin
                valid_6 <= 1'h0;
              end else if (_T_113) begin
                if (4'h6 == idxUnlock_1[3:0]) begin
                  valid_6 <= 1'h0;
                end else begin
                  valid_6 <= _GEN_22;
                end
              end else begin
                valid_6 <= _GEN_22;
              end
            end else if (_T_113) begin
              if (4'h6 == idxUnlock_1[3:0]) begin
                valid_6 <= 1'h0;
              end else begin
                valid_6 <= _GEN_22;
              end
            end else begin
              valid_6 <= _GEN_22;
            end
          end else if (_T_117) begin
            if (4'h6 == idxUnlock_3[3:0]) begin
              valid_6 <= 1'h0;
            end else if (_T_115) begin
              if (4'h6 == idxUnlock_2[3:0]) begin
                valid_6 <= 1'h0;
              end else begin
                valid_6 <= _GEN_54;
              end
            end else begin
              valid_6 <= _GEN_54;
            end
          end else if (_T_115) begin
            if (4'h6 == idxUnlock_2[3:0]) begin
              valid_6 <= 1'h0;
            end else begin
              valid_6 <= _GEN_54;
            end
          end else begin
            valid_6 <= _GEN_54;
          end
        end else if (_T_119) begin
          if (4'h6 == idxUnlock_4[3:0]) begin
            valid_6 <= 1'h0;
          end else if (_T_117) begin
            if (4'h6 == idxUnlock_3[3:0]) begin
              valid_6 <= 1'h0;
            end else begin
              valid_6 <= _GEN_86;
            end
          end else begin
            valid_6 <= _GEN_86;
          end
        end else if (_T_117) begin
          if (4'h6 == idxUnlock_3[3:0]) begin
            valid_6 <= 1'h0;
          end else begin
            valid_6 <= _GEN_86;
          end
        end else begin
          valid_6 <= _GEN_86;
        end
      end else if (_T_121) begin
        if (4'h6 == idxUnlock_5[3:0]) begin
          valid_6 <= 1'h0;
        end else if (_T_119) begin
          if (4'h6 == idxUnlock_4[3:0]) begin
            valid_6 <= 1'h0;
          end else begin
            valid_6 <= _GEN_118;
          end
        end else begin
          valid_6 <= _GEN_118;
        end
      end else if (_T_119) begin
        if (4'h6 == idxUnlock_4[3:0]) begin
          valid_6 <= 1'h0;
        end else begin
          valid_6 <= _GEN_118;
        end
      end else begin
        valid_6 <= _GEN_118;
      end
    end else if (_T_123) begin
      if (4'h6 == idxUnlock_6[3:0]) begin
        valid_6 <= 1'h0;
      end else if (_T_121) begin
        if (4'h6 == idxUnlock_5[3:0]) begin
          valid_6 <= 1'h0;
        end else begin
          valid_6 <= _GEN_150;
        end
      end else begin
        valid_6 <= _GEN_150;
      end
    end else if (_T_121) begin
      if (4'h6 == idxUnlock_5[3:0]) begin
        valid_6 <= 1'h0;
      end else begin
        valid_6 <= _GEN_150;
      end
    end else begin
      valid_6 <= _GEN_150;
    end
    if (reset) begin
      valid_7 <= 1'h0;
    end else if (write) begin
      valid_7 <= _GEN_312;
    end else if (_T_125) begin
      if (4'h7 == idxUnlock_7[3:0]) begin
        valid_7 <= 1'h0;
      end else if (_T_123) begin
        if (4'h7 == idxUnlock_6[3:0]) begin
          valid_7 <= 1'h0;
        end else if (_T_121) begin
          if (4'h7 == idxUnlock_5[3:0]) begin
            valid_7 <= 1'h0;
          end else if (_T_119) begin
            if (4'h7 == idxUnlock_4[3:0]) begin
              valid_7 <= 1'h0;
            end else if (_T_117) begin
              if (4'h7 == idxUnlock_3[3:0]) begin
                valid_7 <= 1'h0;
              end else if (_T_115) begin
                if (4'h7 == idxUnlock_2[3:0]) begin
                  valid_7 <= 1'h0;
                end else if (_T_113) begin
                  if (4'h7 == idxUnlock_1[3:0]) begin
                    valid_7 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'h7 == idxUnlock_0[3:0]) begin
                      valid_7 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h7 == idxUnlock_0[3:0]) begin
                    valid_7 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'h7 == idxUnlock_1[3:0]) begin
                  valid_7 <= 1'h0;
                end else if (_T_111) begin
                  if (4'h7 == idxUnlock_0[3:0]) begin
                    valid_7 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'h7 == idxUnlock_0[3:0]) begin
                  valid_7 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'h7 == idxUnlock_2[3:0]) begin
                valid_7 <= 1'h0;
              end else if (_T_113) begin
                if (4'h7 == idxUnlock_1[3:0]) begin
                  valid_7 <= 1'h0;
                end else begin
                  valid_7 <= _GEN_23;
                end
              end else begin
                valid_7 <= _GEN_23;
              end
            end else if (_T_113) begin
              if (4'h7 == idxUnlock_1[3:0]) begin
                valid_7 <= 1'h0;
              end else begin
                valid_7 <= _GEN_23;
              end
            end else begin
              valid_7 <= _GEN_23;
            end
          end else if (_T_117) begin
            if (4'h7 == idxUnlock_3[3:0]) begin
              valid_7 <= 1'h0;
            end else if (_T_115) begin
              if (4'h7 == idxUnlock_2[3:0]) begin
                valid_7 <= 1'h0;
              end else begin
                valid_7 <= _GEN_55;
              end
            end else begin
              valid_7 <= _GEN_55;
            end
          end else if (_T_115) begin
            if (4'h7 == idxUnlock_2[3:0]) begin
              valid_7 <= 1'h0;
            end else begin
              valid_7 <= _GEN_55;
            end
          end else begin
            valid_7 <= _GEN_55;
          end
        end else if (_T_119) begin
          if (4'h7 == idxUnlock_4[3:0]) begin
            valid_7 <= 1'h0;
          end else if (_T_117) begin
            if (4'h7 == idxUnlock_3[3:0]) begin
              valid_7 <= 1'h0;
            end else begin
              valid_7 <= _GEN_87;
            end
          end else begin
            valid_7 <= _GEN_87;
          end
        end else if (_T_117) begin
          if (4'h7 == idxUnlock_3[3:0]) begin
            valid_7 <= 1'h0;
          end else begin
            valid_7 <= _GEN_87;
          end
        end else begin
          valid_7 <= _GEN_87;
        end
      end else if (_T_121) begin
        if (4'h7 == idxUnlock_5[3:0]) begin
          valid_7 <= 1'h0;
        end else if (_T_119) begin
          if (4'h7 == idxUnlock_4[3:0]) begin
            valid_7 <= 1'h0;
          end else begin
            valid_7 <= _GEN_119;
          end
        end else begin
          valid_7 <= _GEN_119;
        end
      end else if (_T_119) begin
        if (4'h7 == idxUnlock_4[3:0]) begin
          valid_7 <= 1'h0;
        end else begin
          valid_7 <= _GEN_119;
        end
      end else begin
        valid_7 <= _GEN_119;
      end
    end else if (_T_123) begin
      if (4'h7 == idxUnlock_6[3:0]) begin
        valid_7 <= 1'h0;
      end else if (_T_121) begin
        if (4'h7 == idxUnlock_5[3:0]) begin
          valid_7 <= 1'h0;
        end else begin
          valid_7 <= _GEN_151;
        end
      end else begin
        valid_7 <= _GEN_151;
      end
    end else if (_T_121) begin
      if (4'h7 == idxUnlock_5[3:0]) begin
        valid_7 <= 1'h0;
      end else begin
        valid_7 <= _GEN_151;
      end
    end else begin
      valid_7 <= _GEN_151;
    end
    if (reset) begin
      valid_8 <= 1'h0;
    end else if (write) begin
      valid_8 <= _GEN_313;
    end else if (_T_125) begin
      if (4'h8 == idxUnlock_7[3:0]) begin
        valid_8 <= 1'h0;
      end else if (_T_123) begin
        if (4'h8 == idxUnlock_6[3:0]) begin
          valid_8 <= 1'h0;
        end else if (_T_121) begin
          if (4'h8 == idxUnlock_5[3:0]) begin
            valid_8 <= 1'h0;
          end else if (_T_119) begin
            if (4'h8 == idxUnlock_4[3:0]) begin
              valid_8 <= 1'h0;
            end else if (_T_117) begin
              if (4'h8 == idxUnlock_3[3:0]) begin
                valid_8 <= 1'h0;
              end else if (_T_115) begin
                if (4'h8 == idxUnlock_2[3:0]) begin
                  valid_8 <= 1'h0;
                end else if (_T_113) begin
                  if (4'h8 == idxUnlock_1[3:0]) begin
                    valid_8 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'h8 == idxUnlock_0[3:0]) begin
                      valid_8 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h8 == idxUnlock_0[3:0]) begin
                    valid_8 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'h8 == idxUnlock_1[3:0]) begin
                  valid_8 <= 1'h0;
                end else if (_T_111) begin
                  if (4'h8 == idxUnlock_0[3:0]) begin
                    valid_8 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'h8 == idxUnlock_0[3:0]) begin
                  valid_8 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'h8 == idxUnlock_2[3:0]) begin
                valid_8 <= 1'h0;
              end else if (_T_113) begin
                if (4'h8 == idxUnlock_1[3:0]) begin
                  valid_8 <= 1'h0;
                end else begin
                  valid_8 <= _GEN_24;
                end
              end else begin
                valid_8 <= _GEN_24;
              end
            end else if (_T_113) begin
              if (4'h8 == idxUnlock_1[3:0]) begin
                valid_8 <= 1'h0;
              end else begin
                valid_8 <= _GEN_24;
              end
            end else begin
              valid_8 <= _GEN_24;
            end
          end else if (_T_117) begin
            if (4'h8 == idxUnlock_3[3:0]) begin
              valid_8 <= 1'h0;
            end else if (_T_115) begin
              if (4'h8 == idxUnlock_2[3:0]) begin
                valid_8 <= 1'h0;
              end else begin
                valid_8 <= _GEN_56;
              end
            end else begin
              valid_8 <= _GEN_56;
            end
          end else if (_T_115) begin
            if (4'h8 == idxUnlock_2[3:0]) begin
              valid_8 <= 1'h0;
            end else begin
              valid_8 <= _GEN_56;
            end
          end else begin
            valid_8 <= _GEN_56;
          end
        end else if (_T_119) begin
          if (4'h8 == idxUnlock_4[3:0]) begin
            valid_8 <= 1'h0;
          end else if (_T_117) begin
            if (4'h8 == idxUnlock_3[3:0]) begin
              valid_8 <= 1'h0;
            end else begin
              valid_8 <= _GEN_88;
            end
          end else begin
            valid_8 <= _GEN_88;
          end
        end else if (_T_117) begin
          if (4'h8 == idxUnlock_3[3:0]) begin
            valid_8 <= 1'h0;
          end else begin
            valid_8 <= _GEN_88;
          end
        end else begin
          valid_8 <= _GEN_88;
        end
      end else if (_T_121) begin
        if (4'h8 == idxUnlock_5[3:0]) begin
          valid_8 <= 1'h0;
        end else if (_T_119) begin
          if (4'h8 == idxUnlock_4[3:0]) begin
            valid_8 <= 1'h0;
          end else begin
            valid_8 <= _GEN_120;
          end
        end else begin
          valid_8 <= _GEN_120;
        end
      end else if (_T_119) begin
        if (4'h8 == idxUnlock_4[3:0]) begin
          valid_8 <= 1'h0;
        end else begin
          valid_8 <= _GEN_120;
        end
      end else begin
        valid_8 <= _GEN_120;
      end
    end else if (_T_123) begin
      if (4'h8 == idxUnlock_6[3:0]) begin
        valid_8 <= 1'h0;
      end else if (_T_121) begin
        if (4'h8 == idxUnlock_5[3:0]) begin
          valid_8 <= 1'h0;
        end else begin
          valid_8 <= _GEN_152;
        end
      end else begin
        valid_8 <= _GEN_152;
      end
    end else if (_T_121) begin
      if (4'h8 == idxUnlock_5[3:0]) begin
        valid_8 <= 1'h0;
      end else begin
        valid_8 <= _GEN_152;
      end
    end else begin
      valid_8 <= _GEN_152;
    end
    if (reset) begin
      valid_9 <= 1'h0;
    end else if (write) begin
      valid_9 <= _GEN_314;
    end else if (_T_125) begin
      if (4'h9 == idxUnlock_7[3:0]) begin
        valid_9 <= 1'h0;
      end else if (_T_123) begin
        if (4'h9 == idxUnlock_6[3:0]) begin
          valid_9 <= 1'h0;
        end else if (_T_121) begin
          if (4'h9 == idxUnlock_5[3:0]) begin
            valid_9 <= 1'h0;
          end else if (_T_119) begin
            if (4'h9 == idxUnlock_4[3:0]) begin
              valid_9 <= 1'h0;
            end else if (_T_117) begin
              if (4'h9 == idxUnlock_3[3:0]) begin
                valid_9 <= 1'h0;
              end else if (_T_115) begin
                if (4'h9 == idxUnlock_2[3:0]) begin
                  valid_9 <= 1'h0;
                end else if (_T_113) begin
                  if (4'h9 == idxUnlock_1[3:0]) begin
                    valid_9 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'h9 == idxUnlock_0[3:0]) begin
                      valid_9 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'h9 == idxUnlock_0[3:0]) begin
                    valid_9 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'h9 == idxUnlock_1[3:0]) begin
                  valid_9 <= 1'h0;
                end else if (_T_111) begin
                  if (4'h9 == idxUnlock_0[3:0]) begin
                    valid_9 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'h9 == idxUnlock_0[3:0]) begin
                  valid_9 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'h9 == idxUnlock_2[3:0]) begin
                valid_9 <= 1'h0;
              end else if (_T_113) begin
                if (4'h9 == idxUnlock_1[3:0]) begin
                  valid_9 <= 1'h0;
                end else begin
                  valid_9 <= _GEN_25;
                end
              end else begin
                valid_9 <= _GEN_25;
              end
            end else if (_T_113) begin
              if (4'h9 == idxUnlock_1[3:0]) begin
                valid_9 <= 1'h0;
              end else begin
                valid_9 <= _GEN_25;
              end
            end else begin
              valid_9 <= _GEN_25;
            end
          end else if (_T_117) begin
            if (4'h9 == idxUnlock_3[3:0]) begin
              valid_9 <= 1'h0;
            end else if (_T_115) begin
              if (4'h9 == idxUnlock_2[3:0]) begin
                valid_9 <= 1'h0;
              end else begin
                valid_9 <= _GEN_57;
              end
            end else begin
              valid_9 <= _GEN_57;
            end
          end else if (_T_115) begin
            if (4'h9 == idxUnlock_2[3:0]) begin
              valid_9 <= 1'h0;
            end else begin
              valid_9 <= _GEN_57;
            end
          end else begin
            valid_9 <= _GEN_57;
          end
        end else if (_T_119) begin
          if (4'h9 == idxUnlock_4[3:0]) begin
            valid_9 <= 1'h0;
          end else if (_T_117) begin
            if (4'h9 == idxUnlock_3[3:0]) begin
              valid_9 <= 1'h0;
            end else begin
              valid_9 <= _GEN_89;
            end
          end else begin
            valid_9 <= _GEN_89;
          end
        end else if (_T_117) begin
          if (4'h9 == idxUnlock_3[3:0]) begin
            valid_9 <= 1'h0;
          end else begin
            valid_9 <= _GEN_89;
          end
        end else begin
          valid_9 <= _GEN_89;
        end
      end else if (_T_121) begin
        if (4'h9 == idxUnlock_5[3:0]) begin
          valid_9 <= 1'h0;
        end else if (_T_119) begin
          if (4'h9 == idxUnlock_4[3:0]) begin
            valid_9 <= 1'h0;
          end else begin
            valid_9 <= _GEN_121;
          end
        end else begin
          valid_9 <= _GEN_121;
        end
      end else if (_T_119) begin
        if (4'h9 == idxUnlock_4[3:0]) begin
          valid_9 <= 1'h0;
        end else begin
          valid_9 <= _GEN_121;
        end
      end else begin
        valid_9 <= _GEN_121;
      end
    end else if (_T_123) begin
      if (4'h9 == idxUnlock_6[3:0]) begin
        valid_9 <= 1'h0;
      end else if (_T_121) begin
        if (4'h9 == idxUnlock_5[3:0]) begin
          valid_9 <= 1'h0;
        end else begin
          valid_9 <= _GEN_153;
        end
      end else begin
        valid_9 <= _GEN_153;
      end
    end else if (_T_121) begin
      if (4'h9 == idxUnlock_5[3:0]) begin
        valid_9 <= 1'h0;
      end else begin
        valid_9 <= _GEN_153;
      end
    end else begin
      valid_9 <= _GEN_153;
    end
    if (reset) begin
      valid_10 <= 1'h0;
    end else if (write) begin
      valid_10 <= _GEN_315;
    end else if (_T_125) begin
      if (4'ha == idxUnlock_7[3:0]) begin
        valid_10 <= 1'h0;
      end else if (_T_123) begin
        if (4'ha == idxUnlock_6[3:0]) begin
          valid_10 <= 1'h0;
        end else if (_T_121) begin
          if (4'ha == idxUnlock_5[3:0]) begin
            valid_10 <= 1'h0;
          end else if (_T_119) begin
            if (4'ha == idxUnlock_4[3:0]) begin
              valid_10 <= 1'h0;
            end else if (_T_117) begin
              if (4'ha == idxUnlock_3[3:0]) begin
                valid_10 <= 1'h0;
              end else if (_T_115) begin
                if (4'ha == idxUnlock_2[3:0]) begin
                  valid_10 <= 1'h0;
                end else if (_T_113) begin
                  if (4'ha == idxUnlock_1[3:0]) begin
                    valid_10 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'ha == idxUnlock_0[3:0]) begin
                      valid_10 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'ha == idxUnlock_0[3:0]) begin
                    valid_10 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'ha == idxUnlock_1[3:0]) begin
                  valid_10 <= 1'h0;
                end else if (_T_111) begin
                  if (4'ha == idxUnlock_0[3:0]) begin
                    valid_10 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'ha == idxUnlock_0[3:0]) begin
                  valid_10 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'ha == idxUnlock_2[3:0]) begin
                valid_10 <= 1'h0;
              end else if (_T_113) begin
                if (4'ha == idxUnlock_1[3:0]) begin
                  valid_10 <= 1'h0;
                end else begin
                  valid_10 <= _GEN_26;
                end
              end else begin
                valid_10 <= _GEN_26;
              end
            end else if (_T_113) begin
              if (4'ha == idxUnlock_1[3:0]) begin
                valid_10 <= 1'h0;
              end else begin
                valid_10 <= _GEN_26;
              end
            end else begin
              valid_10 <= _GEN_26;
            end
          end else if (_T_117) begin
            if (4'ha == idxUnlock_3[3:0]) begin
              valid_10 <= 1'h0;
            end else if (_T_115) begin
              if (4'ha == idxUnlock_2[3:0]) begin
                valid_10 <= 1'h0;
              end else begin
                valid_10 <= _GEN_58;
              end
            end else begin
              valid_10 <= _GEN_58;
            end
          end else if (_T_115) begin
            if (4'ha == idxUnlock_2[3:0]) begin
              valid_10 <= 1'h0;
            end else begin
              valid_10 <= _GEN_58;
            end
          end else begin
            valid_10 <= _GEN_58;
          end
        end else if (_T_119) begin
          if (4'ha == idxUnlock_4[3:0]) begin
            valid_10 <= 1'h0;
          end else if (_T_117) begin
            if (4'ha == idxUnlock_3[3:0]) begin
              valid_10 <= 1'h0;
            end else begin
              valid_10 <= _GEN_90;
            end
          end else begin
            valid_10 <= _GEN_90;
          end
        end else if (_T_117) begin
          if (4'ha == idxUnlock_3[3:0]) begin
            valid_10 <= 1'h0;
          end else begin
            valid_10 <= _GEN_90;
          end
        end else begin
          valid_10 <= _GEN_90;
        end
      end else if (_T_121) begin
        if (4'ha == idxUnlock_5[3:0]) begin
          valid_10 <= 1'h0;
        end else if (_T_119) begin
          if (4'ha == idxUnlock_4[3:0]) begin
            valid_10 <= 1'h0;
          end else begin
            valid_10 <= _GEN_122;
          end
        end else begin
          valid_10 <= _GEN_122;
        end
      end else if (_T_119) begin
        if (4'ha == idxUnlock_4[3:0]) begin
          valid_10 <= 1'h0;
        end else begin
          valid_10 <= _GEN_122;
        end
      end else begin
        valid_10 <= _GEN_122;
      end
    end else if (_T_123) begin
      if (4'ha == idxUnlock_6[3:0]) begin
        valid_10 <= 1'h0;
      end else if (_T_121) begin
        if (4'ha == idxUnlock_5[3:0]) begin
          valid_10 <= 1'h0;
        end else begin
          valid_10 <= _GEN_154;
        end
      end else begin
        valid_10 <= _GEN_154;
      end
    end else if (_T_121) begin
      if (4'ha == idxUnlock_5[3:0]) begin
        valid_10 <= 1'h0;
      end else begin
        valid_10 <= _GEN_154;
      end
    end else begin
      valid_10 <= _GEN_154;
    end
    if (reset) begin
      valid_11 <= 1'h0;
    end else if (write) begin
      valid_11 <= _GEN_316;
    end else if (_T_125) begin
      if (4'hb == idxUnlock_7[3:0]) begin
        valid_11 <= 1'h0;
      end else if (_T_123) begin
        if (4'hb == idxUnlock_6[3:0]) begin
          valid_11 <= 1'h0;
        end else if (_T_121) begin
          if (4'hb == idxUnlock_5[3:0]) begin
            valid_11 <= 1'h0;
          end else if (_T_119) begin
            if (4'hb == idxUnlock_4[3:0]) begin
              valid_11 <= 1'h0;
            end else if (_T_117) begin
              if (4'hb == idxUnlock_3[3:0]) begin
                valid_11 <= 1'h0;
              end else if (_T_115) begin
                if (4'hb == idxUnlock_2[3:0]) begin
                  valid_11 <= 1'h0;
                end else if (_T_113) begin
                  if (4'hb == idxUnlock_1[3:0]) begin
                    valid_11 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'hb == idxUnlock_0[3:0]) begin
                      valid_11 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'hb == idxUnlock_0[3:0]) begin
                    valid_11 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'hb == idxUnlock_1[3:0]) begin
                  valid_11 <= 1'h0;
                end else if (_T_111) begin
                  if (4'hb == idxUnlock_0[3:0]) begin
                    valid_11 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'hb == idxUnlock_0[3:0]) begin
                  valid_11 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'hb == idxUnlock_2[3:0]) begin
                valid_11 <= 1'h0;
              end else if (_T_113) begin
                if (4'hb == idxUnlock_1[3:0]) begin
                  valid_11 <= 1'h0;
                end else begin
                  valid_11 <= _GEN_27;
                end
              end else begin
                valid_11 <= _GEN_27;
              end
            end else if (_T_113) begin
              if (4'hb == idxUnlock_1[3:0]) begin
                valid_11 <= 1'h0;
              end else begin
                valid_11 <= _GEN_27;
              end
            end else begin
              valid_11 <= _GEN_27;
            end
          end else if (_T_117) begin
            if (4'hb == idxUnlock_3[3:0]) begin
              valid_11 <= 1'h0;
            end else if (_T_115) begin
              if (4'hb == idxUnlock_2[3:0]) begin
                valid_11 <= 1'h0;
              end else begin
                valid_11 <= _GEN_59;
              end
            end else begin
              valid_11 <= _GEN_59;
            end
          end else if (_T_115) begin
            if (4'hb == idxUnlock_2[3:0]) begin
              valid_11 <= 1'h0;
            end else begin
              valid_11 <= _GEN_59;
            end
          end else begin
            valid_11 <= _GEN_59;
          end
        end else if (_T_119) begin
          if (4'hb == idxUnlock_4[3:0]) begin
            valid_11 <= 1'h0;
          end else if (_T_117) begin
            if (4'hb == idxUnlock_3[3:0]) begin
              valid_11 <= 1'h0;
            end else begin
              valid_11 <= _GEN_91;
            end
          end else begin
            valid_11 <= _GEN_91;
          end
        end else if (_T_117) begin
          if (4'hb == idxUnlock_3[3:0]) begin
            valid_11 <= 1'h0;
          end else begin
            valid_11 <= _GEN_91;
          end
        end else begin
          valid_11 <= _GEN_91;
        end
      end else if (_T_121) begin
        if (4'hb == idxUnlock_5[3:0]) begin
          valid_11 <= 1'h0;
        end else if (_T_119) begin
          if (4'hb == idxUnlock_4[3:0]) begin
            valid_11 <= 1'h0;
          end else begin
            valid_11 <= _GEN_123;
          end
        end else begin
          valid_11 <= _GEN_123;
        end
      end else if (_T_119) begin
        if (4'hb == idxUnlock_4[3:0]) begin
          valid_11 <= 1'h0;
        end else begin
          valid_11 <= _GEN_123;
        end
      end else begin
        valid_11 <= _GEN_123;
      end
    end else if (_T_123) begin
      if (4'hb == idxUnlock_6[3:0]) begin
        valid_11 <= 1'h0;
      end else if (_T_121) begin
        if (4'hb == idxUnlock_5[3:0]) begin
          valid_11 <= 1'h0;
        end else begin
          valid_11 <= _GEN_155;
        end
      end else begin
        valid_11 <= _GEN_155;
      end
    end else if (_T_121) begin
      if (4'hb == idxUnlock_5[3:0]) begin
        valid_11 <= 1'h0;
      end else begin
        valid_11 <= _GEN_155;
      end
    end else begin
      valid_11 <= _GEN_155;
    end
    if (reset) begin
      valid_12 <= 1'h0;
    end else if (write) begin
      valid_12 <= _GEN_317;
    end else if (_T_125) begin
      if (4'hc == idxUnlock_7[3:0]) begin
        valid_12 <= 1'h0;
      end else if (_T_123) begin
        if (4'hc == idxUnlock_6[3:0]) begin
          valid_12 <= 1'h0;
        end else if (_T_121) begin
          if (4'hc == idxUnlock_5[3:0]) begin
            valid_12 <= 1'h0;
          end else if (_T_119) begin
            if (4'hc == idxUnlock_4[3:0]) begin
              valid_12 <= 1'h0;
            end else if (_T_117) begin
              if (4'hc == idxUnlock_3[3:0]) begin
                valid_12 <= 1'h0;
              end else if (_T_115) begin
                if (4'hc == idxUnlock_2[3:0]) begin
                  valid_12 <= 1'h0;
                end else if (_T_113) begin
                  if (4'hc == idxUnlock_1[3:0]) begin
                    valid_12 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'hc == idxUnlock_0[3:0]) begin
                      valid_12 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'hc == idxUnlock_0[3:0]) begin
                    valid_12 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'hc == idxUnlock_1[3:0]) begin
                  valid_12 <= 1'h0;
                end else if (_T_111) begin
                  if (4'hc == idxUnlock_0[3:0]) begin
                    valid_12 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'hc == idxUnlock_0[3:0]) begin
                  valid_12 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'hc == idxUnlock_2[3:0]) begin
                valid_12 <= 1'h0;
              end else if (_T_113) begin
                if (4'hc == idxUnlock_1[3:0]) begin
                  valid_12 <= 1'h0;
                end else begin
                  valid_12 <= _GEN_28;
                end
              end else begin
                valid_12 <= _GEN_28;
              end
            end else if (_T_113) begin
              if (4'hc == idxUnlock_1[3:0]) begin
                valid_12 <= 1'h0;
              end else begin
                valid_12 <= _GEN_28;
              end
            end else begin
              valid_12 <= _GEN_28;
            end
          end else if (_T_117) begin
            if (4'hc == idxUnlock_3[3:0]) begin
              valid_12 <= 1'h0;
            end else if (_T_115) begin
              if (4'hc == idxUnlock_2[3:0]) begin
                valid_12 <= 1'h0;
              end else begin
                valid_12 <= _GEN_60;
              end
            end else begin
              valid_12 <= _GEN_60;
            end
          end else if (_T_115) begin
            if (4'hc == idxUnlock_2[3:0]) begin
              valid_12 <= 1'h0;
            end else begin
              valid_12 <= _GEN_60;
            end
          end else begin
            valid_12 <= _GEN_60;
          end
        end else if (_T_119) begin
          if (4'hc == idxUnlock_4[3:0]) begin
            valid_12 <= 1'h0;
          end else if (_T_117) begin
            if (4'hc == idxUnlock_3[3:0]) begin
              valid_12 <= 1'h0;
            end else begin
              valid_12 <= _GEN_92;
            end
          end else begin
            valid_12 <= _GEN_92;
          end
        end else if (_T_117) begin
          if (4'hc == idxUnlock_3[3:0]) begin
            valid_12 <= 1'h0;
          end else begin
            valid_12 <= _GEN_92;
          end
        end else begin
          valid_12 <= _GEN_92;
        end
      end else if (_T_121) begin
        if (4'hc == idxUnlock_5[3:0]) begin
          valid_12 <= 1'h0;
        end else if (_T_119) begin
          if (4'hc == idxUnlock_4[3:0]) begin
            valid_12 <= 1'h0;
          end else begin
            valid_12 <= _GEN_124;
          end
        end else begin
          valid_12 <= _GEN_124;
        end
      end else if (_T_119) begin
        if (4'hc == idxUnlock_4[3:0]) begin
          valid_12 <= 1'h0;
        end else begin
          valid_12 <= _GEN_124;
        end
      end else begin
        valid_12 <= _GEN_124;
      end
    end else if (_T_123) begin
      if (4'hc == idxUnlock_6[3:0]) begin
        valid_12 <= 1'h0;
      end else if (_T_121) begin
        if (4'hc == idxUnlock_5[3:0]) begin
          valid_12 <= 1'h0;
        end else begin
          valid_12 <= _GEN_156;
        end
      end else begin
        valid_12 <= _GEN_156;
      end
    end else if (_T_121) begin
      if (4'hc == idxUnlock_5[3:0]) begin
        valid_12 <= 1'h0;
      end else begin
        valid_12 <= _GEN_156;
      end
    end else begin
      valid_12 <= _GEN_156;
    end
    if (reset) begin
      valid_13 <= 1'h0;
    end else if (write) begin
      valid_13 <= _GEN_318;
    end else if (_T_125) begin
      if (4'hd == idxUnlock_7[3:0]) begin
        valid_13 <= 1'h0;
      end else if (_T_123) begin
        if (4'hd == idxUnlock_6[3:0]) begin
          valid_13 <= 1'h0;
        end else if (_T_121) begin
          if (4'hd == idxUnlock_5[3:0]) begin
            valid_13 <= 1'h0;
          end else if (_T_119) begin
            if (4'hd == idxUnlock_4[3:0]) begin
              valid_13 <= 1'h0;
            end else if (_T_117) begin
              if (4'hd == idxUnlock_3[3:0]) begin
                valid_13 <= 1'h0;
              end else if (_T_115) begin
                if (4'hd == idxUnlock_2[3:0]) begin
                  valid_13 <= 1'h0;
                end else if (_T_113) begin
                  if (4'hd == idxUnlock_1[3:0]) begin
                    valid_13 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'hd == idxUnlock_0[3:0]) begin
                      valid_13 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'hd == idxUnlock_0[3:0]) begin
                    valid_13 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'hd == idxUnlock_1[3:0]) begin
                  valid_13 <= 1'h0;
                end else if (_T_111) begin
                  if (4'hd == idxUnlock_0[3:0]) begin
                    valid_13 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'hd == idxUnlock_0[3:0]) begin
                  valid_13 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'hd == idxUnlock_2[3:0]) begin
                valid_13 <= 1'h0;
              end else if (_T_113) begin
                if (4'hd == idxUnlock_1[3:0]) begin
                  valid_13 <= 1'h0;
                end else begin
                  valid_13 <= _GEN_29;
                end
              end else begin
                valid_13 <= _GEN_29;
              end
            end else if (_T_113) begin
              if (4'hd == idxUnlock_1[3:0]) begin
                valid_13 <= 1'h0;
              end else begin
                valid_13 <= _GEN_29;
              end
            end else begin
              valid_13 <= _GEN_29;
            end
          end else if (_T_117) begin
            if (4'hd == idxUnlock_3[3:0]) begin
              valid_13 <= 1'h0;
            end else if (_T_115) begin
              if (4'hd == idxUnlock_2[3:0]) begin
                valid_13 <= 1'h0;
              end else begin
                valid_13 <= _GEN_61;
              end
            end else begin
              valid_13 <= _GEN_61;
            end
          end else if (_T_115) begin
            if (4'hd == idxUnlock_2[3:0]) begin
              valid_13 <= 1'h0;
            end else begin
              valid_13 <= _GEN_61;
            end
          end else begin
            valid_13 <= _GEN_61;
          end
        end else if (_T_119) begin
          if (4'hd == idxUnlock_4[3:0]) begin
            valid_13 <= 1'h0;
          end else if (_T_117) begin
            if (4'hd == idxUnlock_3[3:0]) begin
              valid_13 <= 1'h0;
            end else begin
              valid_13 <= _GEN_93;
            end
          end else begin
            valid_13 <= _GEN_93;
          end
        end else if (_T_117) begin
          if (4'hd == idxUnlock_3[3:0]) begin
            valid_13 <= 1'h0;
          end else begin
            valid_13 <= _GEN_93;
          end
        end else begin
          valid_13 <= _GEN_93;
        end
      end else if (_T_121) begin
        if (4'hd == idxUnlock_5[3:0]) begin
          valid_13 <= 1'h0;
        end else if (_T_119) begin
          if (4'hd == idxUnlock_4[3:0]) begin
            valid_13 <= 1'h0;
          end else begin
            valid_13 <= _GEN_125;
          end
        end else begin
          valid_13 <= _GEN_125;
        end
      end else if (_T_119) begin
        if (4'hd == idxUnlock_4[3:0]) begin
          valid_13 <= 1'h0;
        end else begin
          valid_13 <= _GEN_125;
        end
      end else begin
        valid_13 <= _GEN_125;
      end
    end else if (_T_123) begin
      if (4'hd == idxUnlock_6[3:0]) begin
        valid_13 <= 1'h0;
      end else if (_T_121) begin
        if (4'hd == idxUnlock_5[3:0]) begin
          valid_13 <= 1'h0;
        end else begin
          valid_13 <= _GEN_157;
        end
      end else begin
        valid_13 <= _GEN_157;
      end
    end else if (_T_121) begin
      if (4'hd == idxUnlock_5[3:0]) begin
        valid_13 <= 1'h0;
      end else begin
        valid_13 <= _GEN_157;
      end
    end else begin
      valid_13 <= _GEN_157;
    end
    if (reset) begin
      valid_14 <= 1'h0;
    end else if (write) begin
      valid_14 <= _GEN_319;
    end else if (_T_125) begin
      if (4'he == idxUnlock_7[3:0]) begin
        valid_14 <= 1'h0;
      end else if (_T_123) begin
        if (4'he == idxUnlock_6[3:0]) begin
          valid_14 <= 1'h0;
        end else if (_T_121) begin
          if (4'he == idxUnlock_5[3:0]) begin
            valid_14 <= 1'h0;
          end else if (_T_119) begin
            if (4'he == idxUnlock_4[3:0]) begin
              valid_14 <= 1'h0;
            end else if (_T_117) begin
              if (4'he == idxUnlock_3[3:0]) begin
                valid_14 <= 1'h0;
              end else if (_T_115) begin
                if (4'he == idxUnlock_2[3:0]) begin
                  valid_14 <= 1'h0;
                end else if (_T_113) begin
                  if (4'he == idxUnlock_1[3:0]) begin
                    valid_14 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'he == idxUnlock_0[3:0]) begin
                      valid_14 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'he == idxUnlock_0[3:0]) begin
                    valid_14 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'he == idxUnlock_1[3:0]) begin
                  valid_14 <= 1'h0;
                end else if (_T_111) begin
                  if (4'he == idxUnlock_0[3:0]) begin
                    valid_14 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'he == idxUnlock_0[3:0]) begin
                  valid_14 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'he == idxUnlock_2[3:0]) begin
                valid_14 <= 1'h0;
              end else if (_T_113) begin
                if (4'he == idxUnlock_1[3:0]) begin
                  valid_14 <= 1'h0;
                end else begin
                  valid_14 <= _GEN_30;
                end
              end else begin
                valid_14 <= _GEN_30;
              end
            end else if (_T_113) begin
              if (4'he == idxUnlock_1[3:0]) begin
                valid_14 <= 1'h0;
              end else begin
                valid_14 <= _GEN_30;
              end
            end else begin
              valid_14 <= _GEN_30;
            end
          end else if (_T_117) begin
            if (4'he == idxUnlock_3[3:0]) begin
              valid_14 <= 1'h0;
            end else if (_T_115) begin
              if (4'he == idxUnlock_2[3:0]) begin
                valid_14 <= 1'h0;
              end else begin
                valid_14 <= _GEN_62;
              end
            end else begin
              valid_14 <= _GEN_62;
            end
          end else if (_T_115) begin
            if (4'he == idxUnlock_2[3:0]) begin
              valid_14 <= 1'h0;
            end else begin
              valid_14 <= _GEN_62;
            end
          end else begin
            valid_14 <= _GEN_62;
          end
        end else if (_T_119) begin
          if (4'he == idxUnlock_4[3:0]) begin
            valid_14 <= 1'h0;
          end else if (_T_117) begin
            if (4'he == idxUnlock_3[3:0]) begin
              valid_14 <= 1'h0;
            end else begin
              valid_14 <= _GEN_94;
            end
          end else begin
            valid_14 <= _GEN_94;
          end
        end else if (_T_117) begin
          if (4'he == idxUnlock_3[3:0]) begin
            valid_14 <= 1'h0;
          end else begin
            valid_14 <= _GEN_94;
          end
        end else begin
          valid_14 <= _GEN_94;
        end
      end else if (_T_121) begin
        if (4'he == idxUnlock_5[3:0]) begin
          valid_14 <= 1'h0;
        end else if (_T_119) begin
          if (4'he == idxUnlock_4[3:0]) begin
            valid_14 <= 1'h0;
          end else begin
            valid_14 <= _GEN_126;
          end
        end else begin
          valid_14 <= _GEN_126;
        end
      end else if (_T_119) begin
        if (4'he == idxUnlock_4[3:0]) begin
          valid_14 <= 1'h0;
        end else begin
          valid_14 <= _GEN_126;
        end
      end else begin
        valid_14 <= _GEN_126;
      end
    end else if (_T_123) begin
      if (4'he == idxUnlock_6[3:0]) begin
        valid_14 <= 1'h0;
      end else if (_T_121) begin
        if (4'he == idxUnlock_5[3:0]) begin
          valid_14 <= 1'h0;
        end else begin
          valid_14 <= _GEN_158;
        end
      end else begin
        valid_14 <= _GEN_158;
      end
    end else if (_T_121) begin
      if (4'he == idxUnlock_5[3:0]) begin
        valid_14 <= 1'h0;
      end else begin
        valid_14 <= _GEN_158;
      end
    end else begin
      valid_14 <= _GEN_158;
    end
    if (reset) begin
      valid_15 <= 1'h0;
    end else if (write) begin
      valid_15 <= _GEN_320;
    end else if (_T_125) begin
      if (4'hf == idxUnlock_7[3:0]) begin
        valid_15 <= 1'h0;
      end else if (_T_123) begin
        if (4'hf == idxUnlock_6[3:0]) begin
          valid_15 <= 1'h0;
        end else if (_T_121) begin
          if (4'hf == idxUnlock_5[3:0]) begin
            valid_15 <= 1'h0;
          end else if (_T_119) begin
            if (4'hf == idxUnlock_4[3:0]) begin
              valid_15 <= 1'h0;
            end else if (_T_117) begin
              if (4'hf == idxUnlock_3[3:0]) begin
                valid_15 <= 1'h0;
              end else if (_T_115) begin
                if (4'hf == idxUnlock_2[3:0]) begin
                  valid_15 <= 1'h0;
                end else if (_T_113) begin
                  if (4'hf == idxUnlock_1[3:0]) begin
                    valid_15 <= 1'h0;
                  end else if (_T_111) begin
                    if (4'hf == idxUnlock_0[3:0]) begin
                      valid_15 <= 1'h0;
                    end
                  end
                end else if (_T_111) begin
                  if (4'hf == idxUnlock_0[3:0]) begin
                    valid_15 <= 1'h0;
                  end
                end
              end else if (_T_113) begin
                if (4'hf == idxUnlock_1[3:0]) begin
                  valid_15 <= 1'h0;
                end else if (_T_111) begin
                  if (4'hf == idxUnlock_0[3:0]) begin
                    valid_15 <= 1'h0;
                  end
                end
              end else if (_T_111) begin
                if (4'hf == idxUnlock_0[3:0]) begin
                  valid_15 <= 1'h0;
                end
              end
            end else if (_T_115) begin
              if (4'hf == idxUnlock_2[3:0]) begin
                valid_15 <= 1'h0;
              end else if (_T_113) begin
                if (4'hf == idxUnlock_1[3:0]) begin
                  valid_15 <= 1'h0;
                end else begin
                  valid_15 <= _GEN_31;
                end
              end else begin
                valid_15 <= _GEN_31;
              end
            end else if (_T_113) begin
              if (4'hf == idxUnlock_1[3:0]) begin
                valid_15 <= 1'h0;
              end else begin
                valid_15 <= _GEN_31;
              end
            end else begin
              valid_15 <= _GEN_31;
            end
          end else if (_T_117) begin
            if (4'hf == idxUnlock_3[3:0]) begin
              valid_15 <= 1'h0;
            end else if (_T_115) begin
              if (4'hf == idxUnlock_2[3:0]) begin
                valid_15 <= 1'h0;
              end else begin
                valid_15 <= _GEN_63;
              end
            end else begin
              valid_15 <= _GEN_63;
            end
          end else if (_T_115) begin
            if (4'hf == idxUnlock_2[3:0]) begin
              valid_15 <= 1'h0;
            end else begin
              valid_15 <= _GEN_63;
            end
          end else begin
            valid_15 <= _GEN_63;
          end
        end else if (_T_119) begin
          if (4'hf == idxUnlock_4[3:0]) begin
            valid_15 <= 1'h0;
          end else if (_T_117) begin
            if (4'hf == idxUnlock_3[3:0]) begin
              valid_15 <= 1'h0;
            end else begin
              valid_15 <= _GEN_95;
            end
          end else begin
            valid_15 <= _GEN_95;
          end
        end else if (_T_117) begin
          if (4'hf == idxUnlock_3[3:0]) begin
            valid_15 <= 1'h0;
          end else begin
            valid_15 <= _GEN_95;
          end
        end else begin
          valid_15 <= _GEN_95;
        end
      end else if (_T_121) begin
        if (4'hf == idxUnlock_5[3:0]) begin
          valid_15 <= 1'h0;
        end else if (_T_119) begin
          if (4'hf == idxUnlock_4[3:0]) begin
            valid_15 <= 1'h0;
          end else begin
            valid_15 <= _GEN_127;
          end
        end else begin
          valid_15 <= _GEN_127;
        end
      end else if (_T_119) begin
        if (4'hf == idxUnlock_4[3:0]) begin
          valid_15 <= 1'h0;
        end else begin
          valid_15 <= _GEN_127;
        end
      end else begin
        valid_15 <= _GEN_127;
      end
    end else if (_T_123) begin
      if (4'hf == idxUnlock_6[3:0]) begin
        valid_15 <= 1'h0;
      end else if (_T_121) begin
        if (4'hf == idxUnlock_5[3:0]) begin
          valid_15 <= 1'h0;
        end else begin
          valid_15 <= _GEN_159;
        end
      end else begin
        valid_15 <= _GEN_159;
      end
    end else if (_T_121) begin
      if (4'hf == idxUnlock_5[3:0]) begin
        valid_15 <= 1'h0;
      end else begin
        valid_15 <= _GEN_159;
      end
    end else begin
      valid_15 <= _GEN_159;
    end
  end
endmodule
module stateMem(
  input         clock,
  input         reset,
  input         io_in_0_valid,
  input  [1:0]  io_in_0_bits_state_state,
  input  [31:0] io_in_0_bits_addr,
  input  [1:0]  io_in_0_bits_way,
  input         io_in_1_valid,
  input  [1:0]  io_in_1_bits_state_state,
  input  [31:0] io_in_1_bits_addr,
  input  [1:0]  io_in_1_bits_way,
  input         io_in_2_valid,
  input  [1:0]  io_in_2_bits_state_state,
  input  [31:0] io_in_2_bits_addr,
  input  [1:0]  io_in_2_bits_way,
  input         io_in_3_valid,
  input  [1:0]  io_in_3_bits_state_state,
  input  [31:0] io_in_3_bits_addr,
  input  [1:0]  io_in_3_bits_way,
  input         io_in_4_valid,
  input  [1:0]  io_in_4_bits_state_state,
  input  [31:0] io_in_4_bits_addr,
  input  [1:0]  io_in_4_bits_way,
  input         io_in_5_valid,
  input  [1:0]  io_in_5_bits_state_state,
  input  [31:0] io_in_5_bits_addr,
  input  [1:0]  io_in_5_bits_way,
  input         io_in_6_valid,
  input  [1:0]  io_in_6_bits_state_state,
  input  [31:0] io_in_6_bits_addr,
  input  [1:0]  io_in_6_bits_way,
  input         io_in_7_valid,
  input  [1:0]  io_in_7_bits_state_state,
  input  [31:0] io_in_7_bits_addr,
  input  [1:0]  io_in_7_bits_way,
  input         io_in_8_valid,
  input  [31:0] io_in_8_bits_addr,
  input  [1:0]  io_in_8_bits_way,
  output        io_out_valid,
  output [1:0]  io_out_bits_state
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] states_0_state; // @[elements.scala 234:25]
  reg [1:0] states_1_state; // @[elements.scala 234:25]
  reg [1:0] states_2_state; // @[elements.scala 234:25]
  reg [1:0] states_3_state; // @[elements.scala 234:25]
  wire  _T_7 = io_in_8_bits_way != 2'h2; // @[elements.scala 237:91]
  wire  isGet = io_in_8_valid & _T_7; // @[elements.scala 237:66]
  wire  _T_9 = io_in_0_bits_way != 2'h2; // @[elements.scala 243:81]
  wire  isSet_0 = io_in_0_valid & _T_9; // @[elements.scala 243:61]
  wire [1:0] _GEN_68 = {{1'd0}, io_in_0_bits_addr[0]}; // @[elements.scala 244:88]
  wire [2:0] _T_13 = _GEN_68 * 2'h2; // @[elements.scala 244:88]
  wire [2:0] _GEN_69 = {{1'd0}, io_in_0_bits_way}; // @[elements.scala 244:98]
  wire [2:0] _T_15 = _T_13 + _GEN_69; // @[elements.scala 244:98]
  wire [2:0] _T_16 = _T_9 ? _T_15 : 3'h0; // @[elements.scala 244:26]
  wire  _T_18 = io_in_1_bits_way != 2'h2; // @[elements.scala 243:81]
  wire  isSet_1 = io_in_1_valid & _T_18; // @[elements.scala 243:61]
  wire [1:0] _GEN_70 = {{1'd0}, io_in_1_bits_addr[0]}; // @[elements.scala 244:88]
  wire [2:0] _T_22 = _GEN_70 * 2'h2; // @[elements.scala 244:88]
  wire [2:0] _GEN_71 = {{1'd0}, io_in_1_bits_way}; // @[elements.scala 244:98]
  wire [2:0] _T_24 = _T_22 + _GEN_71; // @[elements.scala 244:98]
  wire [2:0] _T_25 = _T_18 ? _T_24 : 3'h0; // @[elements.scala 244:26]
  wire  _T_27 = io_in_2_bits_way != 2'h2; // @[elements.scala 243:81]
  wire  isSet_2 = io_in_2_valid & _T_27; // @[elements.scala 243:61]
  wire [1:0] _GEN_72 = {{1'd0}, io_in_2_bits_addr[0]}; // @[elements.scala 244:88]
  wire [2:0] _T_31 = _GEN_72 * 2'h2; // @[elements.scala 244:88]
  wire [2:0] _GEN_73 = {{1'd0}, io_in_2_bits_way}; // @[elements.scala 244:98]
  wire [2:0] _T_33 = _T_31 + _GEN_73; // @[elements.scala 244:98]
  wire [2:0] _T_34 = _T_27 ? _T_33 : 3'h0; // @[elements.scala 244:26]
  wire  _T_36 = io_in_3_bits_way != 2'h2; // @[elements.scala 243:81]
  wire  isSet_3 = io_in_3_valid & _T_36; // @[elements.scala 243:61]
  wire [1:0] _GEN_74 = {{1'd0}, io_in_3_bits_addr[0]}; // @[elements.scala 244:88]
  wire [2:0] _T_40 = _GEN_74 * 2'h2; // @[elements.scala 244:88]
  wire [2:0] _GEN_75 = {{1'd0}, io_in_3_bits_way}; // @[elements.scala 244:98]
  wire [2:0] _T_42 = _T_40 + _GEN_75; // @[elements.scala 244:98]
  wire [2:0] _T_43 = _T_36 ? _T_42 : 3'h0; // @[elements.scala 244:26]
  wire  _T_45 = io_in_4_bits_way != 2'h2; // @[elements.scala 243:81]
  wire  isSet_4 = io_in_4_valid & _T_45; // @[elements.scala 243:61]
  wire [1:0] _GEN_76 = {{1'd0}, io_in_4_bits_addr[0]}; // @[elements.scala 244:88]
  wire [2:0] _T_49 = _GEN_76 * 2'h2; // @[elements.scala 244:88]
  wire [2:0] _GEN_77 = {{1'd0}, io_in_4_bits_way}; // @[elements.scala 244:98]
  wire [2:0] _T_51 = _T_49 + _GEN_77; // @[elements.scala 244:98]
  wire [2:0] _T_52 = _T_45 ? _T_51 : 3'h0; // @[elements.scala 244:26]
  wire  _T_54 = io_in_5_bits_way != 2'h2; // @[elements.scala 243:81]
  wire  isSet_5 = io_in_5_valid & _T_54; // @[elements.scala 243:61]
  wire [1:0] _GEN_78 = {{1'd0}, io_in_5_bits_addr[0]}; // @[elements.scala 244:88]
  wire [2:0] _T_58 = _GEN_78 * 2'h2; // @[elements.scala 244:88]
  wire [2:0] _GEN_79 = {{1'd0}, io_in_5_bits_way}; // @[elements.scala 244:98]
  wire [2:0] _T_60 = _T_58 + _GEN_79; // @[elements.scala 244:98]
  wire [2:0] _T_61 = _T_54 ? _T_60 : 3'h0; // @[elements.scala 244:26]
  wire  _T_63 = io_in_6_bits_way != 2'h2; // @[elements.scala 243:81]
  wire  isSet_6 = io_in_6_valid & _T_63; // @[elements.scala 243:61]
  wire [1:0] _GEN_80 = {{1'd0}, io_in_6_bits_addr[0]}; // @[elements.scala 244:88]
  wire [2:0] _T_67 = _GEN_80 * 2'h2; // @[elements.scala 244:88]
  wire [2:0] _GEN_81 = {{1'd0}, io_in_6_bits_way}; // @[elements.scala 244:98]
  wire [2:0] _T_69 = _T_67 + _GEN_81; // @[elements.scala 244:98]
  wire [2:0] _T_70 = _T_63 ? _T_69 : 3'h0; // @[elements.scala 244:26]
  wire  _T_72 = io_in_7_bits_way != 2'h2; // @[elements.scala 243:81]
  wire  isSet_7 = io_in_7_valid & _T_72; // @[elements.scala 243:61]
  wire [1:0] _GEN_82 = {{1'd0}, io_in_7_bits_addr[0]}; // @[elements.scala 244:88]
  wire [2:0] _T_76 = _GEN_82 * 2'h2; // @[elements.scala 244:88]
  wire [2:0] _GEN_83 = {{1'd0}, io_in_7_bits_way}; // @[elements.scala 244:98]
  wire [2:0] _T_78 = _T_76 + _GEN_83; // @[elements.scala 244:98]
  wire [2:0] _T_79 = _T_72 ? _T_78 : 3'h0; // @[elements.scala 244:26]
  wire [1:0] idxSet_0 = _T_16[1:0]; // @[elements.scala 240:23 elements.scala 244:20]
  wire [1:0] _GEN_0 = 2'h0 == idxSet_0 ? io_in_0_bits_state_state : states_0_state; // @[elements.scala 249:31]
  wire [1:0] _GEN_1 = 2'h1 == idxSet_0 ? io_in_0_bits_state_state : states_1_state; // @[elements.scala 249:31]
  wire [1:0] _GEN_2 = 2'h2 == idxSet_0 ? io_in_0_bits_state_state : states_2_state; // @[elements.scala 249:31]
  wire [1:0] _GEN_3 = 2'h3 == idxSet_0 ? io_in_0_bits_state_state : states_3_state; // @[elements.scala 249:31]
  wire [1:0] _GEN_4 = isSet_0 ? _GEN_0 : states_0_state; // @[elements.scala 248:24]
  wire [1:0] _GEN_5 = isSet_0 ? _GEN_1 : states_1_state; // @[elements.scala 248:24]
  wire [1:0] _GEN_6 = isSet_0 ? _GEN_2 : states_2_state; // @[elements.scala 248:24]
  wire [1:0] _GEN_7 = isSet_0 ? _GEN_3 : states_3_state; // @[elements.scala 248:24]
  wire [1:0] idxSet_1 = _T_25[1:0]; // @[elements.scala 240:23 elements.scala 244:20]
  wire [1:0] _GEN_8 = 2'h0 == idxSet_1 ? io_in_1_bits_state_state : _GEN_4; // @[elements.scala 249:31]
  wire [1:0] _GEN_9 = 2'h1 == idxSet_1 ? io_in_1_bits_state_state : _GEN_5; // @[elements.scala 249:31]
  wire [1:0] _GEN_10 = 2'h2 == idxSet_1 ? io_in_1_bits_state_state : _GEN_6; // @[elements.scala 249:31]
  wire [1:0] _GEN_11 = 2'h3 == idxSet_1 ? io_in_1_bits_state_state : _GEN_7; // @[elements.scala 249:31]
  wire [1:0] _GEN_12 = isSet_1 ? _GEN_8 : _GEN_4; // @[elements.scala 248:24]
  wire [1:0] _GEN_13 = isSet_1 ? _GEN_9 : _GEN_5; // @[elements.scala 248:24]
  wire [1:0] _GEN_14 = isSet_1 ? _GEN_10 : _GEN_6; // @[elements.scala 248:24]
  wire [1:0] _GEN_15 = isSet_1 ? _GEN_11 : _GEN_7; // @[elements.scala 248:24]
  wire [1:0] idxSet_2 = _T_34[1:0]; // @[elements.scala 240:23 elements.scala 244:20]
  wire [1:0] _GEN_16 = 2'h0 == idxSet_2 ? io_in_2_bits_state_state : _GEN_12; // @[elements.scala 249:31]
  wire [1:0] _GEN_17 = 2'h1 == idxSet_2 ? io_in_2_bits_state_state : _GEN_13; // @[elements.scala 249:31]
  wire [1:0] _GEN_18 = 2'h2 == idxSet_2 ? io_in_2_bits_state_state : _GEN_14; // @[elements.scala 249:31]
  wire [1:0] _GEN_19 = 2'h3 == idxSet_2 ? io_in_2_bits_state_state : _GEN_15; // @[elements.scala 249:31]
  wire [1:0] _GEN_20 = isSet_2 ? _GEN_16 : _GEN_12; // @[elements.scala 248:24]
  wire [1:0] _GEN_21 = isSet_2 ? _GEN_17 : _GEN_13; // @[elements.scala 248:24]
  wire [1:0] _GEN_22 = isSet_2 ? _GEN_18 : _GEN_14; // @[elements.scala 248:24]
  wire [1:0] _GEN_23 = isSet_2 ? _GEN_19 : _GEN_15; // @[elements.scala 248:24]
  wire [1:0] idxSet_3 = _T_43[1:0]; // @[elements.scala 240:23 elements.scala 244:20]
  wire [1:0] _GEN_24 = 2'h0 == idxSet_3 ? io_in_3_bits_state_state : _GEN_20; // @[elements.scala 249:31]
  wire [1:0] _GEN_25 = 2'h1 == idxSet_3 ? io_in_3_bits_state_state : _GEN_21; // @[elements.scala 249:31]
  wire [1:0] _GEN_26 = 2'h2 == idxSet_3 ? io_in_3_bits_state_state : _GEN_22; // @[elements.scala 249:31]
  wire [1:0] _GEN_27 = 2'h3 == idxSet_3 ? io_in_3_bits_state_state : _GEN_23; // @[elements.scala 249:31]
  wire [1:0] _GEN_28 = isSet_3 ? _GEN_24 : _GEN_20; // @[elements.scala 248:24]
  wire [1:0] _GEN_29 = isSet_3 ? _GEN_25 : _GEN_21; // @[elements.scala 248:24]
  wire [1:0] _GEN_30 = isSet_3 ? _GEN_26 : _GEN_22; // @[elements.scala 248:24]
  wire [1:0] _GEN_31 = isSet_3 ? _GEN_27 : _GEN_23; // @[elements.scala 248:24]
  wire [1:0] idxSet_4 = _T_52[1:0]; // @[elements.scala 240:23 elements.scala 244:20]
  wire [1:0] _GEN_32 = 2'h0 == idxSet_4 ? io_in_4_bits_state_state : _GEN_28; // @[elements.scala 249:31]
  wire [1:0] _GEN_33 = 2'h1 == idxSet_4 ? io_in_4_bits_state_state : _GEN_29; // @[elements.scala 249:31]
  wire [1:0] _GEN_34 = 2'h2 == idxSet_4 ? io_in_4_bits_state_state : _GEN_30; // @[elements.scala 249:31]
  wire [1:0] _GEN_35 = 2'h3 == idxSet_4 ? io_in_4_bits_state_state : _GEN_31; // @[elements.scala 249:31]
  wire [1:0] _GEN_36 = isSet_4 ? _GEN_32 : _GEN_28; // @[elements.scala 248:24]
  wire [1:0] _GEN_37 = isSet_4 ? _GEN_33 : _GEN_29; // @[elements.scala 248:24]
  wire [1:0] _GEN_38 = isSet_4 ? _GEN_34 : _GEN_30; // @[elements.scala 248:24]
  wire [1:0] _GEN_39 = isSet_4 ? _GEN_35 : _GEN_31; // @[elements.scala 248:24]
  wire [1:0] idxSet_5 = _T_61[1:0]; // @[elements.scala 240:23 elements.scala 244:20]
  wire [1:0] idxSet_6 = _T_70[1:0]; // @[elements.scala 240:23 elements.scala 244:20]
  wire [1:0] idxSet_7 = _T_79[1:0]; // @[elements.scala 240:23 elements.scala 244:20]
  wire [1:0] _GEN_84 = {{1'd0}, io_in_8_bits_addr[0]}; // @[elements.scala 253:91]
  wire [2:0] _T_82 = _GEN_84 * 2'h2; // @[elements.scala 253:91]
  wire [2:0] _GEN_85 = {{1'd0}, io_in_8_bits_way}; // @[elements.scala 253:101]
  wire [2:0] _T_84 = _T_82 + _GEN_85; // @[elements.scala 253:101]
  wire [2:0] _T_85 = _T_7 ? _T_84 : 3'h0; // @[elements.scala 253:19]
  wire [1:0] idxGet = _T_85[1:0]; // @[elements.scala 239:22 elements.scala 253:12]
  wire [1:0] _GEN_65 = 2'h1 == idxGet ? states_1_state : states_0_state; // @[elements.scala 254:17]
  wire [1:0] _GEN_66 = 2'h2 == idxGet ? states_2_state : _GEN_65; // @[elements.scala 254:17]
  assign io_out_valid = _T_7 & isGet; // @[elements.scala 255:18]
  assign io_out_bits_state = 2'h3 == idxGet ? states_3_state : _GEN_66; // @[elements.scala 254:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_0_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  states_1_state = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  states_2_state = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  states_3_state = _RAND_3[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      states_0_state <= 2'h0;
    end else if (isSet_7) begin
      if (2'h0 == idxSet_7) begin
        states_0_state <= io_in_7_bits_state_state;
      end else if (isSet_6) begin
        if (2'h0 == idxSet_6) begin
          states_0_state <= io_in_6_bits_state_state;
        end else if (isSet_5) begin
          if (2'h0 == idxSet_5) begin
            states_0_state <= io_in_5_bits_state_state;
          end else if (isSet_4) begin
            if (2'h0 == idxSet_4) begin
              states_0_state <= io_in_4_bits_state_state;
            end else if (isSet_3) begin
              if (2'h0 == idxSet_3) begin
                states_0_state <= io_in_3_bits_state_state;
              end else if (isSet_2) begin
                if (2'h0 == idxSet_2) begin
                  states_0_state <= io_in_2_bits_state_state;
                end else if (isSet_1) begin
                  if (2'h0 == idxSet_1) begin
                    states_0_state <= io_in_1_bits_state_state;
                  end else if (isSet_0) begin
                    if (2'h0 == idxSet_0) begin
                      states_0_state <= io_in_0_bits_state_state;
                    end
                  end
                end else if (isSet_0) begin
                  if (2'h0 == idxSet_0) begin
                    states_0_state <= io_in_0_bits_state_state;
                  end
                end
              end else if (isSet_1) begin
                if (2'h0 == idxSet_1) begin
                  states_0_state <= io_in_1_bits_state_state;
                end else if (isSet_0) begin
                  if (2'h0 == idxSet_0) begin
                    states_0_state <= io_in_0_bits_state_state;
                  end
                end
              end else if (isSet_0) begin
                if (2'h0 == idxSet_0) begin
                  states_0_state <= io_in_0_bits_state_state;
                end
              end
            end else if (isSet_2) begin
              if (2'h0 == idxSet_2) begin
                states_0_state <= io_in_2_bits_state_state;
              end else if (isSet_1) begin
                if (2'h0 == idxSet_1) begin
                  states_0_state <= io_in_1_bits_state_state;
                end else begin
                  states_0_state <= _GEN_4;
                end
              end else begin
                states_0_state <= _GEN_4;
              end
            end else if (isSet_1) begin
              if (2'h0 == idxSet_1) begin
                states_0_state <= io_in_1_bits_state_state;
              end else begin
                states_0_state <= _GEN_4;
              end
            end else begin
              states_0_state <= _GEN_4;
            end
          end else if (isSet_3) begin
            if (2'h0 == idxSet_3) begin
              states_0_state <= io_in_3_bits_state_state;
            end else if (isSet_2) begin
              if (2'h0 == idxSet_2) begin
                states_0_state <= io_in_2_bits_state_state;
              end else begin
                states_0_state <= _GEN_12;
              end
            end else begin
              states_0_state <= _GEN_12;
            end
          end else if (isSet_2) begin
            if (2'h0 == idxSet_2) begin
              states_0_state <= io_in_2_bits_state_state;
            end else begin
              states_0_state <= _GEN_12;
            end
          end else begin
            states_0_state <= _GEN_12;
          end
        end else if (isSet_4) begin
          if (2'h0 == idxSet_4) begin
            states_0_state <= io_in_4_bits_state_state;
          end else if (isSet_3) begin
            if (2'h0 == idxSet_3) begin
              states_0_state <= io_in_3_bits_state_state;
            end else begin
              states_0_state <= _GEN_20;
            end
          end else begin
            states_0_state <= _GEN_20;
          end
        end else if (isSet_3) begin
          if (2'h0 == idxSet_3) begin
            states_0_state <= io_in_3_bits_state_state;
          end else begin
            states_0_state <= _GEN_20;
          end
        end else begin
          states_0_state <= _GEN_20;
        end
      end else if (isSet_5) begin
        if (2'h0 == idxSet_5) begin
          states_0_state <= io_in_5_bits_state_state;
        end else if (isSet_4) begin
          if (2'h0 == idxSet_4) begin
            states_0_state <= io_in_4_bits_state_state;
          end else begin
            states_0_state <= _GEN_28;
          end
        end else begin
          states_0_state <= _GEN_28;
        end
      end else if (isSet_4) begin
        if (2'h0 == idxSet_4) begin
          states_0_state <= io_in_4_bits_state_state;
        end else begin
          states_0_state <= _GEN_28;
        end
      end else begin
        states_0_state <= _GEN_28;
      end
    end else if (isSet_6) begin
      if (2'h0 == idxSet_6) begin
        states_0_state <= io_in_6_bits_state_state;
      end else if (isSet_5) begin
        if (2'h0 == idxSet_5) begin
          states_0_state <= io_in_5_bits_state_state;
        end else begin
          states_0_state <= _GEN_36;
        end
      end else begin
        states_0_state <= _GEN_36;
      end
    end else if (isSet_5) begin
      if (2'h0 == idxSet_5) begin
        states_0_state <= io_in_5_bits_state_state;
      end else begin
        states_0_state <= _GEN_36;
      end
    end else begin
      states_0_state <= _GEN_36;
    end
    if (reset) begin
      states_1_state <= 2'h0;
    end else if (isSet_7) begin
      if (2'h1 == idxSet_7) begin
        states_1_state <= io_in_7_bits_state_state;
      end else if (isSet_6) begin
        if (2'h1 == idxSet_6) begin
          states_1_state <= io_in_6_bits_state_state;
        end else if (isSet_5) begin
          if (2'h1 == idxSet_5) begin
            states_1_state <= io_in_5_bits_state_state;
          end else if (isSet_4) begin
            if (2'h1 == idxSet_4) begin
              states_1_state <= io_in_4_bits_state_state;
            end else if (isSet_3) begin
              if (2'h1 == idxSet_3) begin
                states_1_state <= io_in_3_bits_state_state;
              end else if (isSet_2) begin
                if (2'h1 == idxSet_2) begin
                  states_1_state <= io_in_2_bits_state_state;
                end else if (isSet_1) begin
                  if (2'h1 == idxSet_1) begin
                    states_1_state <= io_in_1_bits_state_state;
                  end else if (isSet_0) begin
                    if (2'h1 == idxSet_0) begin
                      states_1_state <= io_in_0_bits_state_state;
                    end
                  end
                end else if (isSet_0) begin
                  if (2'h1 == idxSet_0) begin
                    states_1_state <= io_in_0_bits_state_state;
                  end
                end
              end else if (isSet_1) begin
                if (2'h1 == idxSet_1) begin
                  states_1_state <= io_in_1_bits_state_state;
                end else if (isSet_0) begin
                  if (2'h1 == idxSet_0) begin
                    states_1_state <= io_in_0_bits_state_state;
                  end
                end
              end else if (isSet_0) begin
                if (2'h1 == idxSet_0) begin
                  states_1_state <= io_in_0_bits_state_state;
                end
              end
            end else if (isSet_2) begin
              if (2'h1 == idxSet_2) begin
                states_1_state <= io_in_2_bits_state_state;
              end else if (isSet_1) begin
                if (2'h1 == idxSet_1) begin
                  states_1_state <= io_in_1_bits_state_state;
                end else begin
                  states_1_state <= _GEN_5;
                end
              end else begin
                states_1_state <= _GEN_5;
              end
            end else if (isSet_1) begin
              if (2'h1 == idxSet_1) begin
                states_1_state <= io_in_1_bits_state_state;
              end else begin
                states_1_state <= _GEN_5;
              end
            end else begin
              states_1_state <= _GEN_5;
            end
          end else if (isSet_3) begin
            if (2'h1 == idxSet_3) begin
              states_1_state <= io_in_3_bits_state_state;
            end else if (isSet_2) begin
              if (2'h1 == idxSet_2) begin
                states_1_state <= io_in_2_bits_state_state;
              end else begin
                states_1_state <= _GEN_13;
              end
            end else begin
              states_1_state <= _GEN_13;
            end
          end else if (isSet_2) begin
            if (2'h1 == idxSet_2) begin
              states_1_state <= io_in_2_bits_state_state;
            end else begin
              states_1_state <= _GEN_13;
            end
          end else begin
            states_1_state <= _GEN_13;
          end
        end else if (isSet_4) begin
          if (2'h1 == idxSet_4) begin
            states_1_state <= io_in_4_bits_state_state;
          end else if (isSet_3) begin
            if (2'h1 == idxSet_3) begin
              states_1_state <= io_in_3_bits_state_state;
            end else begin
              states_1_state <= _GEN_21;
            end
          end else begin
            states_1_state <= _GEN_21;
          end
        end else if (isSet_3) begin
          if (2'h1 == idxSet_3) begin
            states_1_state <= io_in_3_bits_state_state;
          end else begin
            states_1_state <= _GEN_21;
          end
        end else begin
          states_1_state <= _GEN_21;
        end
      end else if (isSet_5) begin
        if (2'h1 == idxSet_5) begin
          states_1_state <= io_in_5_bits_state_state;
        end else if (isSet_4) begin
          if (2'h1 == idxSet_4) begin
            states_1_state <= io_in_4_bits_state_state;
          end else begin
            states_1_state <= _GEN_29;
          end
        end else begin
          states_1_state <= _GEN_29;
        end
      end else if (isSet_4) begin
        if (2'h1 == idxSet_4) begin
          states_1_state <= io_in_4_bits_state_state;
        end else begin
          states_1_state <= _GEN_29;
        end
      end else begin
        states_1_state <= _GEN_29;
      end
    end else if (isSet_6) begin
      if (2'h1 == idxSet_6) begin
        states_1_state <= io_in_6_bits_state_state;
      end else if (isSet_5) begin
        if (2'h1 == idxSet_5) begin
          states_1_state <= io_in_5_bits_state_state;
        end else begin
          states_1_state <= _GEN_37;
        end
      end else begin
        states_1_state <= _GEN_37;
      end
    end else if (isSet_5) begin
      if (2'h1 == idxSet_5) begin
        states_1_state <= io_in_5_bits_state_state;
      end else begin
        states_1_state <= _GEN_37;
      end
    end else begin
      states_1_state <= _GEN_37;
    end
    if (reset) begin
      states_2_state <= 2'h0;
    end else if (isSet_7) begin
      if (2'h2 == idxSet_7) begin
        states_2_state <= io_in_7_bits_state_state;
      end else if (isSet_6) begin
        if (2'h2 == idxSet_6) begin
          states_2_state <= io_in_6_bits_state_state;
        end else if (isSet_5) begin
          if (2'h2 == idxSet_5) begin
            states_2_state <= io_in_5_bits_state_state;
          end else if (isSet_4) begin
            if (2'h2 == idxSet_4) begin
              states_2_state <= io_in_4_bits_state_state;
            end else if (isSet_3) begin
              if (2'h2 == idxSet_3) begin
                states_2_state <= io_in_3_bits_state_state;
              end else if (isSet_2) begin
                if (2'h2 == idxSet_2) begin
                  states_2_state <= io_in_2_bits_state_state;
                end else if (isSet_1) begin
                  if (2'h2 == idxSet_1) begin
                    states_2_state <= io_in_1_bits_state_state;
                  end else if (isSet_0) begin
                    if (2'h2 == idxSet_0) begin
                      states_2_state <= io_in_0_bits_state_state;
                    end
                  end
                end else if (isSet_0) begin
                  if (2'h2 == idxSet_0) begin
                    states_2_state <= io_in_0_bits_state_state;
                  end
                end
              end else if (isSet_1) begin
                if (2'h2 == idxSet_1) begin
                  states_2_state <= io_in_1_bits_state_state;
                end else if (isSet_0) begin
                  if (2'h2 == idxSet_0) begin
                    states_2_state <= io_in_0_bits_state_state;
                  end
                end
              end else if (isSet_0) begin
                if (2'h2 == idxSet_0) begin
                  states_2_state <= io_in_0_bits_state_state;
                end
              end
            end else if (isSet_2) begin
              if (2'h2 == idxSet_2) begin
                states_2_state <= io_in_2_bits_state_state;
              end else if (isSet_1) begin
                if (2'h2 == idxSet_1) begin
                  states_2_state <= io_in_1_bits_state_state;
                end else begin
                  states_2_state <= _GEN_6;
                end
              end else begin
                states_2_state <= _GEN_6;
              end
            end else if (isSet_1) begin
              if (2'h2 == idxSet_1) begin
                states_2_state <= io_in_1_bits_state_state;
              end else begin
                states_2_state <= _GEN_6;
              end
            end else begin
              states_2_state <= _GEN_6;
            end
          end else if (isSet_3) begin
            if (2'h2 == idxSet_3) begin
              states_2_state <= io_in_3_bits_state_state;
            end else if (isSet_2) begin
              if (2'h2 == idxSet_2) begin
                states_2_state <= io_in_2_bits_state_state;
              end else begin
                states_2_state <= _GEN_14;
              end
            end else begin
              states_2_state <= _GEN_14;
            end
          end else if (isSet_2) begin
            if (2'h2 == idxSet_2) begin
              states_2_state <= io_in_2_bits_state_state;
            end else begin
              states_2_state <= _GEN_14;
            end
          end else begin
            states_2_state <= _GEN_14;
          end
        end else if (isSet_4) begin
          if (2'h2 == idxSet_4) begin
            states_2_state <= io_in_4_bits_state_state;
          end else if (isSet_3) begin
            if (2'h2 == idxSet_3) begin
              states_2_state <= io_in_3_bits_state_state;
            end else begin
              states_2_state <= _GEN_22;
            end
          end else begin
            states_2_state <= _GEN_22;
          end
        end else if (isSet_3) begin
          if (2'h2 == idxSet_3) begin
            states_2_state <= io_in_3_bits_state_state;
          end else begin
            states_2_state <= _GEN_22;
          end
        end else begin
          states_2_state <= _GEN_22;
        end
      end else if (isSet_5) begin
        if (2'h2 == idxSet_5) begin
          states_2_state <= io_in_5_bits_state_state;
        end else if (isSet_4) begin
          if (2'h2 == idxSet_4) begin
            states_2_state <= io_in_4_bits_state_state;
          end else begin
            states_2_state <= _GEN_30;
          end
        end else begin
          states_2_state <= _GEN_30;
        end
      end else if (isSet_4) begin
        if (2'h2 == idxSet_4) begin
          states_2_state <= io_in_4_bits_state_state;
        end else begin
          states_2_state <= _GEN_30;
        end
      end else begin
        states_2_state <= _GEN_30;
      end
    end else if (isSet_6) begin
      if (2'h2 == idxSet_6) begin
        states_2_state <= io_in_6_bits_state_state;
      end else if (isSet_5) begin
        if (2'h2 == idxSet_5) begin
          states_2_state <= io_in_5_bits_state_state;
        end else begin
          states_2_state <= _GEN_38;
        end
      end else begin
        states_2_state <= _GEN_38;
      end
    end else if (isSet_5) begin
      if (2'h2 == idxSet_5) begin
        states_2_state <= io_in_5_bits_state_state;
      end else begin
        states_2_state <= _GEN_38;
      end
    end else begin
      states_2_state <= _GEN_38;
    end
    if (reset) begin
      states_3_state <= 2'h0;
    end else if (isSet_7) begin
      if (2'h3 == idxSet_7) begin
        states_3_state <= io_in_7_bits_state_state;
      end else if (isSet_6) begin
        if (2'h3 == idxSet_6) begin
          states_3_state <= io_in_6_bits_state_state;
        end else if (isSet_5) begin
          if (2'h3 == idxSet_5) begin
            states_3_state <= io_in_5_bits_state_state;
          end else if (isSet_4) begin
            if (2'h3 == idxSet_4) begin
              states_3_state <= io_in_4_bits_state_state;
            end else if (isSet_3) begin
              if (2'h3 == idxSet_3) begin
                states_3_state <= io_in_3_bits_state_state;
              end else if (isSet_2) begin
                if (2'h3 == idxSet_2) begin
                  states_3_state <= io_in_2_bits_state_state;
                end else if (isSet_1) begin
                  if (2'h3 == idxSet_1) begin
                    states_3_state <= io_in_1_bits_state_state;
                  end else if (isSet_0) begin
                    if (2'h3 == idxSet_0) begin
                      states_3_state <= io_in_0_bits_state_state;
                    end
                  end
                end else if (isSet_0) begin
                  if (2'h3 == idxSet_0) begin
                    states_3_state <= io_in_0_bits_state_state;
                  end
                end
              end else if (isSet_1) begin
                if (2'h3 == idxSet_1) begin
                  states_3_state <= io_in_1_bits_state_state;
                end else if (isSet_0) begin
                  if (2'h3 == idxSet_0) begin
                    states_3_state <= io_in_0_bits_state_state;
                  end
                end
              end else if (isSet_0) begin
                if (2'h3 == idxSet_0) begin
                  states_3_state <= io_in_0_bits_state_state;
                end
              end
            end else if (isSet_2) begin
              if (2'h3 == idxSet_2) begin
                states_3_state <= io_in_2_bits_state_state;
              end else if (isSet_1) begin
                if (2'h3 == idxSet_1) begin
                  states_3_state <= io_in_1_bits_state_state;
                end else begin
                  states_3_state <= _GEN_7;
                end
              end else begin
                states_3_state <= _GEN_7;
              end
            end else if (isSet_1) begin
              if (2'h3 == idxSet_1) begin
                states_3_state <= io_in_1_bits_state_state;
              end else begin
                states_3_state <= _GEN_7;
              end
            end else begin
              states_3_state <= _GEN_7;
            end
          end else if (isSet_3) begin
            if (2'h3 == idxSet_3) begin
              states_3_state <= io_in_3_bits_state_state;
            end else if (isSet_2) begin
              if (2'h3 == idxSet_2) begin
                states_3_state <= io_in_2_bits_state_state;
              end else begin
                states_3_state <= _GEN_15;
              end
            end else begin
              states_3_state <= _GEN_15;
            end
          end else if (isSet_2) begin
            if (2'h3 == idxSet_2) begin
              states_3_state <= io_in_2_bits_state_state;
            end else begin
              states_3_state <= _GEN_15;
            end
          end else begin
            states_3_state <= _GEN_15;
          end
        end else if (isSet_4) begin
          if (2'h3 == idxSet_4) begin
            states_3_state <= io_in_4_bits_state_state;
          end else if (isSet_3) begin
            if (2'h3 == idxSet_3) begin
              states_3_state <= io_in_3_bits_state_state;
            end else begin
              states_3_state <= _GEN_23;
            end
          end else begin
            states_3_state <= _GEN_23;
          end
        end else if (isSet_3) begin
          if (2'h3 == idxSet_3) begin
            states_3_state <= io_in_3_bits_state_state;
          end else begin
            states_3_state <= _GEN_23;
          end
        end else begin
          states_3_state <= _GEN_23;
        end
      end else if (isSet_5) begin
        if (2'h3 == idxSet_5) begin
          states_3_state <= io_in_5_bits_state_state;
        end else if (isSet_4) begin
          if (2'h3 == idxSet_4) begin
            states_3_state <= io_in_4_bits_state_state;
          end else begin
            states_3_state <= _GEN_31;
          end
        end else begin
          states_3_state <= _GEN_31;
        end
      end else if (isSet_4) begin
        if (2'h3 == idxSet_4) begin
          states_3_state <= io_in_4_bits_state_state;
        end else begin
          states_3_state <= _GEN_31;
        end
      end else begin
        states_3_state <= _GEN_31;
      end
    end else if (isSet_6) begin
      if (2'h3 == idxSet_6) begin
        states_3_state <= io_in_6_bits_state_state;
      end else if (isSet_5) begin
        if (2'h3 == idxSet_5) begin
          states_3_state <= io_in_5_bits_state_state;
        end else begin
          states_3_state <= _GEN_39;
        end
      end else begin
        states_3_state <= _GEN_39;
      end
    end else if (isSet_5) begin
      if (2'h3 == idxSet_5) begin
        states_3_state <= io_in_5_bits_state_state;
      end else begin
        states_3_state <= _GEN_39;
      end
    end else begin
      states_3_state <= _GEN_39;
    end
  end
endmodule
module FindEmptyLine_10(
  input        io_data_0,
  input        io_data_1,
  input        io_data_2,
  input        io_data_3,
  input        io_data_4,
  input        io_data_5,
  input        io_data_6,
  input        io_data_7,
  output       io_value_valid,
  output [3:0] io_value_bits
);
  wire  _T = ~io_data_0; // @[elements.scala 74:53]
  wire  _T_1 = ~io_data_1; // @[elements.scala 74:53]
  wire  _T_2 = ~io_data_2; // @[elements.scala 74:53]
  wire  _T_3 = ~io_data_3; // @[elements.scala 74:53]
  wire  _T_4 = ~io_data_4; // @[elements.scala 74:53]
  wire  _T_5 = ~io_data_5; // @[elements.scala 74:53]
  wire  _T_6 = ~io_data_6; // @[elements.scala 74:53]
  wire  _T_7 = ~io_data_7; // @[elements.scala 74:53]
  wire [4:0] _GEN_0 = _T_7 ? 5'h7 : 5'h8; // @[elements.scala 74:66]
  wire [4:0] _GEN_2 = _T_6 ? 5'h6 : _GEN_0; // @[elements.scala 74:66]
  wire  _GEN_3 = _T_6 | _T_7; // @[elements.scala 74:66]
  wire [4:0] _GEN_4 = _T_5 ? 5'h5 : _GEN_2; // @[elements.scala 74:66]
  wire  _GEN_5 = _T_5 | _GEN_3; // @[elements.scala 74:66]
  wire [4:0] _GEN_6 = _T_4 ? 5'h4 : _GEN_4; // @[elements.scala 74:66]
  wire  _GEN_7 = _T_4 | _GEN_5; // @[elements.scala 74:66]
  wire [4:0] _GEN_8 = _T_3 ? 5'h3 : _GEN_6; // @[elements.scala 74:66]
  wire  _GEN_9 = _T_3 | _GEN_7; // @[elements.scala 74:66]
  wire [4:0] _GEN_10 = _T_2 ? 5'h2 : _GEN_8; // @[elements.scala 74:66]
  wire  _GEN_11 = _T_2 | _GEN_9; // @[elements.scala 74:66]
  wire [4:0] _GEN_12 = _T_1 ? 5'h1 : _GEN_10; // @[elements.scala 74:66]
  wire  _GEN_13 = _T_1 | _GEN_11; // @[elements.scala 74:66]
  wire [4:0] idx = _T ? 5'h0 : _GEN_12; // @[elements.scala 74:66]
  assign io_value_valid = _T | _GEN_13; // @[elements.scala 68:20 elements.scala 76:32 elements.scala 76:32 elements.scala 76:32 elements.scala 76:32 elements.scala 76:32 elements.scala 76:32 elements.scala 76:32 elements.scala 76:32]
  assign io_value_bits = idx[3:0]; // @[elements.scala 79:19]
endmodule
module PC(
  input         clock,
  input         reset,
  output        io_write_ready,
  input         io_write_valid,
  input  [31:0] io_write_bits_addr,
  input  [1:0]  io_write_bits_way,
  input  [63:0] io_write_bits_data,
  input  [1:0]  io_write_bits_replaceWay,
  input  [31:0] io_write_bits_tbeFields_0,
  input  [15:0] io_write_bits_pc,
  input  [1:0]  io_read_0_in_bits_data_way,
  input  [15:0] io_read_0_in_bits_data_pc,
  input         io_read_0_in_bits_data_valid,
  output [31:0] io_read_0_out_bits_addr,
  output [1:0]  io_read_0_out_bits_way,
  output [63:0] io_read_0_out_bits_data,
  output [1:0]  io_read_0_out_bits_replaceWay,
  output [31:0] io_read_0_out_bits_tbeFields_0,
  output [15:0] io_read_0_out_bits_pc,
  output        io_read_0_out_bits_valid,
  input  [1:0]  io_read_1_in_bits_data_way,
  input  [15:0] io_read_1_in_bits_data_pc,
  input         io_read_1_in_bits_data_valid,
  output [31:0] io_read_1_out_bits_addr,
  output [1:0]  io_read_1_out_bits_way,
  output [63:0] io_read_1_out_bits_data,
  output [1:0]  io_read_1_out_bits_replaceWay,
  output [31:0] io_read_1_out_bits_tbeFields_0,
  output [15:0] io_read_1_out_bits_pc,
  output        io_read_1_out_bits_valid,
  input  [1:0]  io_read_2_in_bits_data_way,
  input  [15:0] io_read_2_in_bits_data_pc,
  input         io_read_2_in_bits_data_valid,
  output [31:0] io_read_2_out_bits_addr,
  output [1:0]  io_read_2_out_bits_way,
  output [63:0] io_read_2_out_bits_data,
  output [1:0]  io_read_2_out_bits_replaceWay,
  output [31:0] io_read_2_out_bits_tbeFields_0,
  output [15:0] io_read_2_out_bits_pc,
  output        io_read_2_out_bits_valid,
  input  [1:0]  io_read_3_in_bits_data_way,
  input  [15:0] io_read_3_in_bits_data_pc,
  input         io_read_3_in_bits_data_valid,
  output [31:0] io_read_3_out_bits_addr,
  output [1:0]  io_read_3_out_bits_way,
  output [63:0] io_read_3_out_bits_data,
  output [1:0]  io_read_3_out_bits_replaceWay,
  output [31:0] io_read_3_out_bits_tbeFields_0,
  output [15:0] io_read_3_out_bits_pc,
  output        io_read_3_out_bits_valid,
  input  [1:0]  io_read_4_in_bits_data_way,
  input  [15:0] io_read_4_in_bits_data_pc,
  input         io_read_4_in_bits_data_valid,
  output [31:0] io_read_4_out_bits_addr,
  output [1:0]  io_read_4_out_bits_way,
  output [63:0] io_read_4_out_bits_data,
  output [1:0]  io_read_4_out_bits_replaceWay,
  output [31:0] io_read_4_out_bits_tbeFields_0,
  output [15:0] io_read_4_out_bits_pc,
  output        io_read_4_out_bits_valid,
  input  [1:0]  io_read_5_in_bits_data_way,
  input  [15:0] io_read_5_in_bits_data_pc,
  input         io_read_5_in_bits_data_valid,
  output [31:0] io_read_5_out_bits_addr,
  output [1:0]  io_read_5_out_bits_way,
  output [63:0] io_read_5_out_bits_data,
  output [1:0]  io_read_5_out_bits_replaceWay,
  output [31:0] io_read_5_out_bits_tbeFields_0,
  output [15:0] io_read_5_out_bits_pc,
  output        io_read_5_out_bits_valid,
  input  [1:0]  io_read_6_in_bits_data_way,
  input  [15:0] io_read_6_in_bits_data_pc,
  input         io_read_6_in_bits_data_valid,
  output [31:0] io_read_6_out_bits_addr,
  output [1:0]  io_read_6_out_bits_way,
  output [63:0] io_read_6_out_bits_data,
  output [1:0]  io_read_6_out_bits_replaceWay,
  output [31:0] io_read_6_out_bits_tbeFields_0,
  output [15:0] io_read_6_out_bits_pc,
  output        io_read_6_out_bits_valid,
  input  [1:0]  io_read_7_in_bits_data_way,
  input  [15:0] io_read_7_in_bits_data_pc,
  input         io_read_7_in_bits_data_valid,
  output [31:0] io_read_7_out_bits_addr,
  output [1:0]  io_read_7_out_bits_way,
  output [63:0] io_read_7_out_bits_data,
  output [1:0]  io_read_7_out_bits_replaceWay,
  output [31:0] io_read_7_out_bits_tbeFields_0,
  output [15:0] io_read_7_out_bits_pc,
  output        io_read_7_out_bits_valid,
  output        io_isFull
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
`endif // RANDOMIZE_REG_INIT
  wire  findNewLine_io_data_0; // @[elements.scala 278:29]
  wire  findNewLine_io_data_1; // @[elements.scala 278:29]
  wire  findNewLine_io_data_2; // @[elements.scala 278:29]
  wire  findNewLine_io_data_3; // @[elements.scala 278:29]
  wire  findNewLine_io_data_4; // @[elements.scala 278:29]
  wire  findNewLine_io_data_5; // @[elements.scala 278:29]
  wire  findNewLine_io_data_6; // @[elements.scala 278:29]
  wire  findNewLine_io_data_7; // @[elements.scala 278:29]
  wire  findNewLine_io_value_valid; // @[elements.scala 278:29]
  wire [3:0] findNewLine_io_value_bits; // @[elements.scala 278:29]
  reg [31:0] pcContent_0_addr; // @[elements.scala 274:29]
  reg [1:0] pcContent_0_way; // @[elements.scala 274:29]
  reg [63:0] pcContent_0_data; // @[elements.scala 274:29]
  reg [1:0] pcContent_0_replaceWay; // @[elements.scala 274:29]
  reg [31:0] pcContent_0_tbeFields_0; // @[elements.scala 274:29]
  reg [15:0] pcContent_0_pc; // @[elements.scala 274:29]
  reg  pcContent_0_valid; // @[elements.scala 274:29]
  reg [31:0] pcContent_1_addr; // @[elements.scala 274:29]
  reg [1:0] pcContent_1_way; // @[elements.scala 274:29]
  reg [63:0] pcContent_1_data; // @[elements.scala 274:29]
  reg [1:0] pcContent_1_replaceWay; // @[elements.scala 274:29]
  reg [31:0] pcContent_1_tbeFields_0; // @[elements.scala 274:29]
  reg [15:0] pcContent_1_pc; // @[elements.scala 274:29]
  reg  pcContent_1_valid; // @[elements.scala 274:29]
  reg [31:0] pcContent_2_addr; // @[elements.scala 274:29]
  reg [1:0] pcContent_2_way; // @[elements.scala 274:29]
  reg [63:0] pcContent_2_data; // @[elements.scala 274:29]
  reg [1:0] pcContent_2_replaceWay; // @[elements.scala 274:29]
  reg [31:0] pcContent_2_tbeFields_0; // @[elements.scala 274:29]
  reg [15:0] pcContent_2_pc; // @[elements.scala 274:29]
  reg  pcContent_2_valid; // @[elements.scala 274:29]
  reg [31:0] pcContent_3_addr; // @[elements.scala 274:29]
  reg [1:0] pcContent_3_way; // @[elements.scala 274:29]
  reg [63:0] pcContent_3_data; // @[elements.scala 274:29]
  reg [1:0] pcContent_3_replaceWay; // @[elements.scala 274:29]
  reg [31:0] pcContent_3_tbeFields_0; // @[elements.scala 274:29]
  reg [15:0] pcContent_3_pc; // @[elements.scala 274:29]
  reg  pcContent_3_valid; // @[elements.scala 274:29]
  reg [31:0] pcContent_4_addr; // @[elements.scala 274:29]
  reg [1:0] pcContent_4_way; // @[elements.scala 274:29]
  reg [63:0] pcContent_4_data; // @[elements.scala 274:29]
  reg [1:0] pcContent_4_replaceWay; // @[elements.scala 274:29]
  reg [31:0] pcContent_4_tbeFields_0; // @[elements.scala 274:29]
  reg [15:0] pcContent_4_pc; // @[elements.scala 274:29]
  reg  pcContent_4_valid; // @[elements.scala 274:29]
  reg [31:0] pcContent_5_addr; // @[elements.scala 274:29]
  reg [1:0] pcContent_5_way; // @[elements.scala 274:29]
  reg [63:0] pcContent_5_data; // @[elements.scala 274:29]
  reg [1:0] pcContent_5_replaceWay; // @[elements.scala 274:29]
  reg [31:0] pcContent_5_tbeFields_0; // @[elements.scala 274:29]
  reg [15:0] pcContent_5_pc; // @[elements.scala 274:29]
  reg  pcContent_5_valid; // @[elements.scala 274:29]
  reg [31:0] pcContent_6_addr; // @[elements.scala 274:29]
  reg [1:0] pcContent_6_way; // @[elements.scala 274:29]
  reg [63:0] pcContent_6_data; // @[elements.scala 274:29]
  reg [1:0] pcContent_6_replaceWay; // @[elements.scala 274:29]
  reg [31:0] pcContent_6_tbeFields_0; // @[elements.scala 274:29]
  reg [15:0] pcContent_6_pc; // @[elements.scala 274:29]
  reg  pcContent_6_valid; // @[elements.scala 274:29]
  reg [31:0] pcContent_7_addr; // @[elements.scala 274:29]
  reg [1:0] pcContent_7_way; // @[elements.scala 274:29]
  reg [63:0] pcContent_7_data; // @[elements.scala 274:29]
  reg [1:0] pcContent_7_replaceWay; // @[elements.scala 274:29]
  reg [31:0] pcContent_7_tbeFields_0; // @[elements.scala 274:29]
  reg [15:0] pcContent_7_pc; // @[elements.scala 274:29]
  reg  pcContent_7_valid; // @[elements.scala 274:29]
  wire  write = io_write_ready & io_write_valid; // @[Decoupled.scala 40:37]
  wire  _T_316 = ~write; // @[elements.scala 288:14]
  wire [3:0] writeIdx = findNewLine_io_value_bits;
  wire  _T_317 = writeIdx != 4'h0; // @[elements.scala 288:41]
  wire  _T_318 = write & _T_317; // @[elements.scala 288:30]
  wire  _T_319 = _T_316 | _T_318; // @[elements.scala 288:21]
  wire  _GEN_1 = _T_319 ? io_read_0_in_bits_data_valid : pcContent_0_valid; // @[elements.scala 288:50]
  wire  _T_321 = writeIdx != 4'h1; // @[elements.scala 288:41]
  wire  _T_322 = write & _T_321; // @[elements.scala 288:30]
  wire  _T_323 = _T_316 | _T_322; // @[elements.scala 288:21]
  wire  _GEN_4 = _T_323 ? io_read_1_in_bits_data_valid : pcContent_1_valid; // @[elements.scala 288:50]
  wire  _T_325 = writeIdx != 4'h2; // @[elements.scala 288:41]
  wire  _T_326 = write & _T_325; // @[elements.scala 288:30]
  wire  _T_327 = _T_316 | _T_326; // @[elements.scala 288:21]
  wire  _GEN_7 = _T_327 ? io_read_2_in_bits_data_valid : pcContent_2_valid; // @[elements.scala 288:50]
  wire  _T_329 = writeIdx != 4'h3; // @[elements.scala 288:41]
  wire  _T_330 = write & _T_329; // @[elements.scala 288:30]
  wire  _T_331 = _T_316 | _T_330; // @[elements.scala 288:21]
  wire  _GEN_10 = _T_331 ? io_read_3_in_bits_data_valid : pcContent_3_valid; // @[elements.scala 288:50]
  wire  _T_333 = writeIdx != 4'h4; // @[elements.scala 288:41]
  wire  _T_334 = write & _T_333; // @[elements.scala 288:30]
  wire  _T_335 = _T_316 | _T_334; // @[elements.scala 288:21]
  wire  _GEN_13 = _T_335 ? io_read_4_in_bits_data_valid : pcContent_4_valid; // @[elements.scala 288:50]
  wire  _T_337 = writeIdx != 4'h5; // @[elements.scala 288:41]
  wire  _T_338 = write & _T_337; // @[elements.scala 288:30]
  wire  _T_339 = _T_316 | _T_338; // @[elements.scala 288:21]
  wire  _GEN_16 = _T_339 ? io_read_5_in_bits_data_valid : pcContent_5_valid; // @[elements.scala 288:50]
  wire  _T_341 = writeIdx != 4'h6; // @[elements.scala 288:41]
  wire  _T_342 = write & _T_341; // @[elements.scala 288:30]
  wire  _T_343 = _T_316 | _T_342; // @[elements.scala 288:21]
  wire  _GEN_19 = _T_343 ? io_read_6_in_bits_data_valid : pcContent_6_valid; // @[elements.scala 288:50]
  wire  _T_345 = writeIdx != 4'h7; // @[elements.scala 288:41]
  wire  _T_346 = write & _T_345; // @[elements.scala 288:30]
  wire  _T_347 = _T_316 | _T_346; // @[elements.scala 288:21]
  wire  _GEN_22 = _T_347 ? io_read_7_in_bits_data_valid : pcContent_7_valid; // @[elements.scala 288:50]
  wire  _GEN_152 = 3'h0 == writeIdx[2:0]; // @[elements.scala 296:28]
  wire  _GEN_80 = _GEN_152 | _GEN_1; // @[elements.scala 296:28]
  wire  _GEN_153 = 3'h1 == writeIdx[2:0]; // @[elements.scala 296:28]
  wire  _GEN_81 = _GEN_153 | _GEN_4; // @[elements.scala 296:28]
  wire  _GEN_154 = 3'h2 == writeIdx[2:0]; // @[elements.scala 296:28]
  wire  _GEN_82 = _GEN_154 | _GEN_7; // @[elements.scala 296:28]
  wire  _GEN_155 = 3'h3 == writeIdx[2:0]; // @[elements.scala 296:28]
  wire  _GEN_83 = _GEN_155 | _GEN_10; // @[elements.scala 296:28]
  wire  _GEN_156 = 3'h4 == writeIdx[2:0]; // @[elements.scala 296:28]
  wire  _GEN_84 = _GEN_156 | _GEN_13; // @[elements.scala 296:28]
  wire  _GEN_157 = 3'h5 == writeIdx[2:0]; // @[elements.scala 296:28]
  wire  _GEN_85 = _GEN_157 | _GEN_16; // @[elements.scala 296:28]
  wire  _GEN_158 = 3'h6 == writeIdx[2:0]; // @[elements.scala 296:28]
  wire  _GEN_86 = _GEN_158 | _GEN_19; // @[elements.scala 296:28]
  wire  _GEN_159 = 3'h7 == writeIdx[2:0]; // @[elements.scala 296:28]
  wire  _GEN_87 = _GEN_159 | _GEN_22; // @[elements.scala 296:28]
  FindEmptyLine_10 findNewLine ( // @[elements.scala 278:29]
    .io_data_0(findNewLine_io_data_0),
    .io_data_1(findNewLine_io_data_1),
    .io_data_2(findNewLine_io_data_2),
    .io_data_3(findNewLine_io_data_3),
    .io_data_4(findNewLine_io_data_4),
    .io_data_5(findNewLine_io_data_5),
    .io_data_6(findNewLine_io_data_6),
    .io_data_7(findNewLine_io_data_7),
    .io_value_valid(findNewLine_io_value_valid),
    .io_value_bits(findNewLine_io_value_bits)
  );
  assign io_write_ready = findNewLine_io_value_valid; // @[elements.scala 299:20]
  assign io_read_0_out_bits_addr = pcContent_0_addr; // @[elements.scala 283:30]
  assign io_read_0_out_bits_way = pcContent_0_way; // @[elements.scala 283:30]
  assign io_read_0_out_bits_data = pcContent_0_data; // @[elements.scala 283:30]
  assign io_read_0_out_bits_replaceWay = pcContent_0_replaceWay; // @[elements.scala 283:30]
  assign io_read_0_out_bits_tbeFields_0 = pcContent_0_tbeFields_0; // @[elements.scala 283:30]
  assign io_read_0_out_bits_pc = pcContent_0_pc; // @[elements.scala 283:30]
  assign io_read_0_out_bits_valid = pcContent_0_valid; // @[elements.scala 283:30]
  assign io_read_1_out_bits_addr = pcContent_1_addr; // @[elements.scala 283:30]
  assign io_read_1_out_bits_way = pcContent_1_way; // @[elements.scala 283:30]
  assign io_read_1_out_bits_data = pcContent_1_data; // @[elements.scala 283:30]
  assign io_read_1_out_bits_replaceWay = pcContent_1_replaceWay; // @[elements.scala 283:30]
  assign io_read_1_out_bits_tbeFields_0 = pcContent_1_tbeFields_0; // @[elements.scala 283:30]
  assign io_read_1_out_bits_pc = pcContent_1_pc; // @[elements.scala 283:30]
  assign io_read_1_out_bits_valid = pcContent_1_valid; // @[elements.scala 283:30]
  assign io_read_2_out_bits_addr = pcContent_2_addr; // @[elements.scala 283:30]
  assign io_read_2_out_bits_way = pcContent_2_way; // @[elements.scala 283:30]
  assign io_read_2_out_bits_data = pcContent_2_data; // @[elements.scala 283:30]
  assign io_read_2_out_bits_replaceWay = pcContent_2_replaceWay; // @[elements.scala 283:30]
  assign io_read_2_out_bits_tbeFields_0 = pcContent_2_tbeFields_0; // @[elements.scala 283:30]
  assign io_read_2_out_bits_pc = pcContent_2_pc; // @[elements.scala 283:30]
  assign io_read_2_out_bits_valid = pcContent_2_valid; // @[elements.scala 283:30]
  assign io_read_3_out_bits_addr = pcContent_3_addr; // @[elements.scala 283:30]
  assign io_read_3_out_bits_way = pcContent_3_way; // @[elements.scala 283:30]
  assign io_read_3_out_bits_data = pcContent_3_data; // @[elements.scala 283:30]
  assign io_read_3_out_bits_replaceWay = pcContent_3_replaceWay; // @[elements.scala 283:30]
  assign io_read_3_out_bits_tbeFields_0 = pcContent_3_tbeFields_0; // @[elements.scala 283:30]
  assign io_read_3_out_bits_pc = pcContent_3_pc; // @[elements.scala 283:30]
  assign io_read_3_out_bits_valid = pcContent_3_valid; // @[elements.scala 283:30]
  assign io_read_4_out_bits_addr = pcContent_4_addr; // @[elements.scala 283:30]
  assign io_read_4_out_bits_way = pcContent_4_way; // @[elements.scala 283:30]
  assign io_read_4_out_bits_data = pcContent_4_data; // @[elements.scala 283:30]
  assign io_read_4_out_bits_replaceWay = pcContent_4_replaceWay; // @[elements.scala 283:30]
  assign io_read_4_out_bits_tbeFields_0 = pcContent_4_tbeFields_0; // @[elements.scala 283:30]
  assign io_read_4_out_bits_pc = pcContent_4_pc; // @[elements.scala 283:30]
  assign io_read_4_out_bits_valid = pcContent_4_valid; // @[elements.scala 283:30]
  assign io_read_5_out_bits_addr = pcContent_5_addr; // @[elements.scala 283:30]
  assign io_read_5_out_bits_way = pcContent_5_way; // @[elements.scala 283:30]
  assign io_read_5_out_bits_data = pcContent_5_data; // @[elements.scala 283:30]
  assign io_read_5_out_bits_replaceWay = pcContent_5_replaceWay; // @[elements.scala 283:30]
  assign io_read_5_out_bits_tbeFields_0 = pcContent_5_tbeFields_0; // @[elements.scala 283:30]
  assign io_read_5_out_bits_pc = pcContent_5_pc; // @[elements.scala 283:30]
  assign io_read_5_out_bits_valid = pcContent_5_valid; // @[elements.scala 283:30]
  assign io_read_6_out_bits_addr = pcContent_6_addr; // @[elements.scala 283:30]
  assign io_read_6_out_bits_way = pcContent_6_way; // @[elements.scala 283:30]
  assign io_read_6_out_bits_data = pcContent_6_data; // @[elements.scala 283:30]
  assign io_read_6_out_bits_replaceWay = pcContent_6_replaceWay; // @[elements.scala 283:30]
  assign io_read_6_out_bits_tbeFields_0 = pcContent_6_tbeFields_0; // @[elements.scala 283:30]
  assign io_read_6_out_bits_pc = pcContent_6_pc; // @[elements.scala 283:30]
  assign io_read_6_out_bits_valid = pcContent_6_valid; // @[elements.scala 283:30]
  assign io_read_7_out_bits_addr = pcContent_7_addr; // @[elements.scala 283:30]
  assign io_read_7_out_bits_way = pcContent_7_way; // @[elements.scala 283:30]
  assign io_read_7_out_bits_data = pcContent_7_data; // @[elements.scala 283:30]
  assign io_read_7_out_bits_replaceWay = pcContent_7_replaceWay; // @[elements.scala 283:30]
  assign io_read_7_out_bits_tbeFields_0 = pcContent_7_tbeFields_0; // @[elements.scala 283:30]
  assign io_read_7_out_bits_pc = pcContent_7_pc; // @[elements.scala 283:30]
  assign io_read_7_out_bits_valid = pcContent_7_valid; // @[elements.scala 283:30]
  assign io_isFull = ~io_write_ready; // @[elements.scala 300:15]
  assign findNewLine_io_data_0 = pcContent_0_valid; // @[elements.scala 279:25]
  assign findNewLine_io_data_1 = pcContent_1_valid; // @[elements.scala 279:25]
  assign findNewLine_io_data_2 = pcContent_2_valid; // @[elements.scala 279:25]
  assign findNewLine_io_data_3 = pcContent_3_valid; // @[elements.scala 279:25]
  assign findNewLine_io_data_4 = pcContent_4_valid; // @[elements.scala 279:25]
  assign findNewLine_io_data_5 = pcContent_5_valid; // @[elements.scala 279:25]
  assign findNewLine_io_data_6 = pcContent_6_valid; // @[elements.scala 279:25]
  assign findNewLine_io_data_7 = pcContent_7_valid; // @[elements.scala 279:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pcContent_0_addr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  pcContent_0_way = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  pcContent_0_data = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  pcContent_0_replaceWay = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  pcContent_0_tbeFields_0 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  pcContent_0_pc = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  pcContent_0_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pcContent_1_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  pcContent_1_way = _RAND_8[1:0];
  _RAND_9 = {2{`RANDOM}};
  pcContent_1_data = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  pcContent_1_replaceWay = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  pcContent_1_tbeFields_0 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  pcContent_1_pc = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  pcContent_1_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  pcContent_2_addr = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  pcContent_2_way = _RAND_15[1:0];
  _RAND_16 = {2{`RANDOM}};
  pcContent_2_data = _RAND_16[63:0];
  _RAND_17 = {1{`RANDOM}};
  pcContent_2_replaceWay = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  pcContent_2_tbeFields_0 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  pcContent_2_pc = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  pcContent_2_valid = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  pcContent_3_addr = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  pcContent_3_way = _RAND_22[1:0];
  _RAND_23 = {2{`RANDOM}};
  pcContent_3_data = _RAND_23[63:0];
  _RAND_24 = {1{`RANDOM}};
  pcContent_3_replaceWay = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  pcContent_3_tbeFields_0 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  pcContent_3_pc = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  pcContent_3_valid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  pcContent_4_addr = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  pcContent_4_way = _RAND_29[1:0];
  _RAND_30 = {2{`RANDOM}};
  pcContent_4_data = _RAND_30[63:0];
  _RAND_31 = {1{`RANDOM}};
  pcContent_4_replaceWay = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  pcContent_4_tbeFields_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  pcContent_4_pc = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  pcContent_4_valid = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  pcContent_5_addr = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  pcContent_5_way = _RAND_36[1:0];
  _RAND_37 = {2{`RANDOM}};
  pcContent_5_data = _RAND_37[63:0];
  _RAND_38 = {1{`RANDOM}};
  pcContent_5_replaceWay = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  pcContent_5_tbeFields_0 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  pcContent_5_pc = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  pcContent_5_valid = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  pcContent_6_addr = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  pcContent_6_way = _RAND_43[1:0];
  _RAND_44 = {2{`RANDOM}};
  pcContent_6_data = _RAND_44[63:0];
  _RAND_45 = {1{`RANDOM}};
  pcContent_6_replaceWay = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  pcContent_6_tbeFields_0 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  pcContent_6_pc = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  pcContent_6_valid = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  pcContent_7_addr = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  pcContent_7_way = _RAND_50[1:0];
  _RAND_51 = {2{`RANDOM}};
  pcContent_7_data = _RAND_51[63:0];
  _RAND_52 = {1{`RANDOM}};
  pcContent_7_replaceWay = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  pcContent_7_tbeFields_0 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  pcContent_7_pc = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  pcContent_7_valid = _RAND_55[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pcContent_0_addr <= 32'h0;
    end else if (write) begin
      if (3'h0 == writeIdx[2:0]) begin
        pcContent_0_addr <= io_write_bits_addr;
      end
    end
    if (reset) begin
      pcContent_0_way <= 2'h2;
    end else if (write) begin
      if (3'h0 == writeIdx[2:0]) begin
        pcContent_0_way <= io_write_bits_way;
      end else if (_T_319) begin
        pcContent_0_way <= io_read_0_in_bits_data_way;
      end
    end else if (_T_319) begin
      pcContent_0_way <= io_read_0_in_bits_data_way;
    end
    if (reset) begin
      pcContent_0_data <= 64'h0;
    end else if (write) begin
      if (3'h0 == writeIdx[2:0]) begin
        pcContent_0_data <= io_write_bits_data;
      end
    end
    if (reset) begin
      pcContent_0_replaceWay <= 2'h0;
    end else if (write) begin
      if (3'h0 == writeIdx[2:0]) begin
        pcContent_0_replaceWay <= io_write_bits_replaceWay;
      end
    end
    if (reset) begin
      pcContent_0_tbeFields_0 <= 32'h0;
    end else if (write) begin
      if (3'h0 == writeIdx[2:0]) begin
        pcContent_0_tbeFields_0 <= io_write_bits_tbeFields_0;
      end
    end
    if (reset) begin
      pcContent_0_pc <= 16'h0;
    end else if (write) begin
      if (3'h0 == writeIdx[2:0]) begin
        pcContent_0_pc <= io_write_bits_pc;
      end else if (_T_319) begin
        pcContent_0_pc <= io_read_0_in_bits_data_pc;
      end
    end else if (_T_319) begin
      pcContent_0_pc <= io_read_0_in_bits_data_pc;
    end
    if (reset) begin
      pcContent_0_valid <= 1'h0;
    end else if (write) begin
      pcContent_0_valid <= _GEN_80;
    end else if (_T_319) begin
      pcContent_0_valid <= io_read_0_in_bits_data_valid;
    end
    if (reset) begin
      pcContent_1_addr <= 32'h0;
    end else if (write) begin
      if (3'h1 == writeIdx[2:0]) begin
        pcContent_1_addr <= io_write_bits_addr;
      end
    end
    if (reset) begin
      pcContent_1_way <= 2'h2;
    end else if (write) begin
      if (3'h1 == writeIdx[2:0]) begin
        pcContent_1_way <= io_write_bits_way;
      end else if (_T_323) begin
        pcContent_1_way <= io_read_1_in_bits_data_way;
      end
    end else if (_T_323) begin
      pcContent_1_way <= io_read_1_in_bits_data_way;
    end
    if (reset) begin
      pcContent_1_data <= 64'h0;
    end else if (write) begin
      if (3'h1 == writeIdx[2:0]) begin
        pcContent_1_data <= io_write_bits_data;
      end
    end
    if (reset) begin
      pcContent_1_replaceWay <= 2'h0;
    end else if (write) begin
      if (3'h1 == writeIdx[2:0]) begin
        pcContent_1_replaceWay <= io_write_bits_replaceWay;
      end
    end
    if (reset) begin
      pcContent_1_tbeFields_0 <= 32'h0;
    end else if (write) begin
      if (3'h1 == writeIdx[2:0]) begin
        pcContent_1_tbeFields_0 <= io_write_bits_tbeFields_0;
      end
    end
    if (reset) begin
      pcContent_1_pc <= 16'h0;
    end else if (write) begin
      if (3'h1 == writeIdx[2:0]) begin
        pcContent_1_pc <= io_write_bits_pc;
      end else if (_T_323) begin
        pcContent_1_pc <= io_read_1_in_bits_data_pc;
      end
    end else if (_T_323) begin
      pcContent_1_pc <= io_read_1_in_bits_data_pc;
    end
    if (reset) begin
      pcContent_1_valid <= 1'h0;
    end else if (write) begin
      pcContent_1_valid <= _GEN_81;
    end else if (_T_323) begin
      pcContent_1_valid <= io_read_1_in_bits_data_valid;
    end
    if (reset) begin
      pcContent_2_addr <= 32'h0;
    end else if (write) begin
      if (3'h2 == writeIdx[2:0]) begin
        pcContent_2_addr <= io_write_bits_addr;
      end
    end
    if (reset) begin
      pcContent_2_way <= 2'h2;
    end else if (write) begin
      if (3'h2 == writeIdx[2:0]) begin
        pcContent_2_way <= io_write_bits_way;
      end else if (_T_327) begin
        pcContent_2_way <= io_read_2_in_bits_data_way;
      end
    end else if (_T_327) begin
      pcContent_2_way <= io_read_2_in_bits_data_way;
    end
    if (reset) begin
      pcContent_2_data <= 64'h0;
    end else if (write) begin
      if (3'h2 == writeIdx[2:0]) begin
        pcContent_2_data <= io_write_bits_data;
      end
    end
    if (reset) begin
      pcContent_2_replaceWay <= 2'h0;
    end else if (write) begin
      if (3'h2 == writeIdx[2:0]) begin
        pcContent_2_replaceWay <= io_write_bits_replaceWay;
      end
    end
    if (reset) begin
      pcContent_2_tbeFields_0 <= 32'h0;
    end else if (write) begin
      if (3'h2 == writeIdx[2:0]) begin
        pcContent_2_tbeFields_0 <= io_write_bits_tbeFields_0;
      end
    end
    if (reset) begin
      pcContent_2_pc <= 16'h0;
    end else if (write) begin
      if (3'h2 == writeIdx[2:0]) begin
        pcContent_2_pc <= io_write_bits_pc;
      end else if (_T_327) begin
        pcContent_2_pc <= io_read_2_in_bits_data_pc;
      end
    end else if (_T_327) begin
      pcContent_2_pc <= io_read_2_in_bits_data_pc;
    end
    if (reset) begin
      pcContent_2_valid <= 1'h0;
    end else if (write) begin
      pcContent_2_valid <= _GEN_82;
    end else if (_T_327) begin
      pcContent_2_valid <= io_read_2_in_bits_data_valid;
    end
    if (reset) begin
      pcContent_3_addr <= 32'h0;
    end else if (write) begin
      if (3'h3 == writeIdx[2:0]) begin
        pcContent_3_addr <= io_write_bits_addr;
      end
    end
    if (reset) begin
      pcContent_3_way <= 2'h2;
    end else if (write) begin
      if (3'h3 == writeIdx[2:0]) begin
        pcContent_3_way <= io_write_bits_way;
      end else if (_T_331) begin
        pcContent_3_way <= io_read_3_in_bits_data_way;
      end
    end else if (_T_331) begin
      pcContent_3_way <= io_read_3_in_bits_data_way;
    end
    if (reset) begin
      pcContent_3_data <= 64'h0;
    end else if (write) begin
      if (3'h3 == writeIdx[2:0]) begin
        pcContent_3_data <= io_write_bits_data;
      end
    end
    if (reset) begin
      pcContent_3_replaceWay <= 2'h0;
    end else if (write) begin
      if (3'h3 == writeIdx[2:0]) begin
        pcContent_3_replaceWay <= io_write_bits_replaceWay;
      end
    end
    if (reset) begin
      pcContent_3_tbeFields_0 <= 32'h0;
    end else if (write) begin
      if (3'h3 == writeIdx[2:0]) begin
        pcContent_3_tbeFields_0 <= io_write_bits_tbeFields_0;
      end
    end
    if (reset) begin
      pcContent_3_pc <= 16'h0;
    end else if (write) begin
      if (3'h3 == writeIdx[2:0]) begin
        pcContent_3_pc <= io_write_bits_pc;
      end else if (_T_331) begin
        pcContent_3_pc <= io_read_3_in_bits_data_pc;
      end
    end else if (_T_331) begin
      pcContent_3_pc <= io_read_3_in_bits_data_pc;
    end
    if (reset) begin
      pcContent_3_valid <= 1'h0;
    end else if (write) begin
      pcContent_3_valid <= _GEN_83;
    end else if (_T_331) begin
      pcContent_3_valid <= io_read_3_in_bits_data_valid;
    end
    if (reset) begin
      pcContent_4_addr <= 32'h0;
    end else if (write) begin
      if (3'h4 == writeIdx[2:0]) begin
        pcContent_4_addr <= io_write_bits_addr;
      end
    end
    if (reset) begin
      pcContent_4_way <= 2'h2;
    end else if (write) begin
      if (3'h4 == writeIdx[2:0]) begin
        pcContent_4_way <= io_write_bits_way;
      end else if (_T_335) begin
        pcContent_4_way <= io_read_4_in_bits_data_way;
      end
    end else if (_T_335) begin
      pcContent_4_way <= io_read_4_in_bits_data_way;
    end
    if (reset) begin
      pcContent_4_data <= 64'h0;
    end else if (write) begin
      if (3'h4 == writeIdx[2:0]) begin
        pcContent_4_data <= io_write_bits_data;
      end
    end
    if (reset) begin
      pcContent_4_replaceWay <= 2'h0;
    end else if (write) begin
      if (3'h4 == writeIdx[2:0]) begin
        pcContent_4_replaceWay <= io_write_bits_replaceWay;
      end
    end
    if (reset) begin
      pcContent_4_tbeFields_0 <= 32'h0;
    end else if (write) begin
      if (3'h4 == writeIdx[2:0]) begin
        pcContent_4_tbeFields_0 <= io_write_bits_tbeFields_0;
      end
    end
    if (reset) begin
      pcContent_4_pc <= 16'h0;
    end else if (write) begin
      if (3'h4 == writeIdx[2:0]) begin
        pcContent_4_pc <= io_write_bits_pc;
      end else if (_T_335) begin
        pcContent_4_pc <= io_read_4_in_bits_data_pc;
      end
    end else if (_T_335) begin
      pcContent_4_pc <= io_read_4_in_bits_data_pc;
    end
    if (reset) begin
      pcContent_4_valid <= 1'h0;
    end else if (write) begin
      pcContent_4_valid <= _GEN_84;
    end else if (_T_335) begin
      pcContent_4_valid <= io_read_4_in_bits_data_valid;
    end
    if (reset) begin
      pcContent_5_addr <= 32'h0;
    end else if (write) begin
      if (3'h5 == writeIdx[2:0]) begin
        pcContent_5_addr <= io_write_bits_addr;
      end
    end
    if (reset) begin
      pcContent_5_way <= 2'h2;
    end else if (write) begin
      if (3'h5 == writeIdx[2:0]) begin
        pcContent_5_way <= io_write_bits_way;
      end else if (_T_339) begin
        pcContent_5_way <= io_read_5_in_bits_data_way;
      end
    end else if (_T_339) begin
      pcContent_5_way <= io_read_5_in_bits_data_way;
    end
    if (reset) begin
      pcContent_5_data <= 64'h0;
    end else if (write) begin
      if (3'h5 == writeIdx[2:0]) begin
        pcContent_5_data <= io_write_bits_data;
      end
    end
    if (reset) begin
      pcContent_5_replaceWay <= 2'h0;
    end else if (write) begin
      if (3'h5 == writeIdx[2:0]) begin
        pcContent_5_replaceWay <= io_write_bits_replaceWay;
      end
    end
    if (reset) begin
      pcContent_5_tbeFields_0 <= 32'h0;
    end else if (write) begin
      if (3'h5 == writeIdx[2:0]) begin
        pcContent_5_tbeFields_0 <= io_write_bits_tbeFields_0;
      end
    end
    if (reset) begin
      pcContent_5_pc <= 16'h0;
    end else if (write) begin
      if (3'h5 == writeIdx[2:0]) begin
        pcContent_5_pc <= io_write_bits_pc;
      end else if (_T_339) begin
        pcContent_5_pc <= io_read_5_in_bits_data_pc;
      end
    end else if (_T_339) begin
      pcContent_5_pc <= io_read_5_in_bits_data_pc;
    end
    if (reset) begin
      pcContent_5_valid <= 1'h0;
    end else if (write) begin
      pcContent_5_valid <= _GEN_85;
    end else if (_T_339) begin
      pcContent_5_valid <= io_read_5_in_bits_data_valid;
    end
    if (reset) begin
      pcContent_6_addr <= 32'h0;
    end else if (write) begin
      if (3'h6 == writeIdx[2:0]) begin
        pcContent_6_addr <= io_write_bits_addr;
      end
    end
    if (reset) begin
      pcContent_6_way <= 2'h2;
    end else if (write) begin
      if (3'h6 == writeIdx[2:0]) begin
        pcContent_6_way <= io_write_bits_way;
      end else if (_T_343) begin
        pcContent_6_way <= io_read_6_in_bits_data_way;
      end
    end else if (_T_343) begin
      pcContent_6_way <= io_read_6_in_bits_data_way;
    end
    if (reset) begin
      pcContent_6_data <= 64'h0;
    end else if (write) begin
      if (3'h6 == writeIdx[2:0]) begin
        pcContent_6_data <= io_write_bits_data;
      end
    end
    if (reset) begin
      pcContent_6_replaceWay <= 2'h0;
    end else if (write) begin
      if (3'h6 == writeIdx[2:0]) begin
        pcContent_6_replaceWay <= io_write_bits_replaceWay;
      end
    end
    if (reset) begin
      pcContent_6_tbeFields_0 <= 32'h0;
    end else if (write) begin
      if (3'h6 == writeIdx[2:0]) begin
        pcContent_6_tbeFields_0 <= io_write_bits_tbeFields_0;
      end
    end
    if (reset) begin
      pcContent_6_pc <= 16'h0;
    end else if (write) begin
      if (3'h6 == writeIdx[2:0]) begin
        pcContent_6_pc <= io_write_bits_pc;
      end else if (_T_343) begin
        pcContent_6_pc <= io_read_6_in_bits_data_pc;
      end
    end else if (_T_343) begin
      pcContent_6_pc <= io_read_6_in_bits_data_pc;
    end
    if (reset) begin
      pcContent_6_valid <= 1'h0;
    end else if (write) begin
      pcContent_6_valid <= _GEN_86;
    end else if (_T_343) begin
      pcContent_6_valid <= io_read_6_in_bits_data_valid;
    end
    if (reset) begin
      pcContent_7_addr <= 32'h0;
    end else if (write) begin
      if (3'h7 == writeIdx[2:0]) begin
        pcContent_7_addr <= io_write_bits_addr;
      end
    end
    if (reset) begin
      pcContent_7_way <= 2'h2;
    end else if (write) begin
      if (3'h7 == writeIdx[2:0]) begin
        pcContent_7_way <= io_write_bits_way;
      end else if (_T_347) begin
        pcContent_7_way <= io_read_7_in_bits_data_way;
      end
    end else if (_T_347) begin
      pcContent_7_way <= io_read_7_in_bits_data_way;
    end
    if (reset) begin
      pcContent_7_data <= 64'h0;
    end else if (write) begin
      if (3'h7 == writeIdx[2:0]) begin
        pcContent_7_data <= io_write_bits_data;
      end
    end
    if (reset) begin
      pcContent_7_replaceWay <= 2'h0;
    end else if (write) begin
      if (3'h7 == writeIdx[2:0]) begin
        pcContent_7_replaceWay <= io_write_bits_replaceWay;
      end
    end
    if (reset) begin
      pcContent_7_tbeFields_0 <= 32'h0;
    end else if (write) begin
      if (3'h7 == writeIdx[2:0]) begin
        pcContent_7_tbeFields_0 <= io_write_bits_tbeFields_0;
      end
    end
    if (reset) begin
      pcContent_7_pc <= 16'h0;
    end else if (write) begin
      if (3'h7 == writeIdx[2:0]) begin
        pcContent_7_pc <= io_write_bits_pc;
      end else if (_T_347) begin
        pcContent_7_pc <= io_read_7_in_bits_data_pc;
      end
    end else if (_T_347) begin
      pcContent_7_pc <= io_read_7_in_bits_data_pc;
    end
    if (reset) begin
      pcContent_7_valid <= 1'h0;
    end else if (write) begin
      pcContent_7_valid <= _GEN_87;
    end else if (_T_347) begin
      pcContent_7_valid <= io_read_7_in_bits_data_valid;
    end
  end
endmodule
module Arbiter_3(
  input         io_in_0_valid,
  input  [1:0]  io_in_0_bits_event,
  input  [31:0] io_in_0_bits_addr,
  input  [63:0] io_in_0_bits_data,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [1:0]  io_in_1_bits_event,
  input  [31:0] io_in_1_bits_addr,
  input  [63:0] io_in_1_bits_data,
  input         io_in_2_valid,
  input  [1:0]  io_in_2_bits_event,
  input  [31:0] io_in_2_bits_addr,
  input  [63:0] io_in_2_bits_data,
  input         io_in_3_valid,
  input  [1:0]  io_in_3_bits_event,
  input  [31:0] io_in_3_bits_addr,
  input  [63:0] io_in_3_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output [1:0]  io_out_bits_event,
  output [31:0] io_out_bits_addr,
  output [63:0] io_out_bits_data,
  output [1:0]  io_chosen
);
  wire [1:0] _GEN_0 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_1 = io_in_2_valid ? io_in_2_bits_data : io_in_3_bits_data; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_2 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_3 = io_in_2_valid ? io_in_2_bits_event : io_in_3_bits_event; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_4 = io_in_1_valid ? 2'h1 : _GEN_0; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_5 = io_in_1_valid ? io_in_1_bits_data : _GEN_1; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_6 = io_in_1_valid ? io_in_1_bits_addr : _GEN_2; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_7 = io_in_1_valid ? io_in_1_bits_event : _GEN_3; // @[Arbiter.scala 126:27]
  wire  _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  _T_1 = _T | io_in_2_valid; // @[Arbiter.scala 31:68]
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  grant_3 = ~_T_1; // @[Arbiter.scala 31:78]
  wire  _T_6 = ~grant_3; // @[Arbiter.scala 135:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_6 | io_in_3_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_event = io_in_0_valid ? io_in_0_bits_event : _GEN_7; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_6; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : _GEN_5; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_chosen = io_in_0_valid ? 2'h0 : _GEN_4; // @[Arbiter.scala 123:13 Arbiter.scala 127:17 Arbiter.scala 127:17 Arbiter.scala 127:17]
endmodule
module RRArbiter_2(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_req_addr,
  input  [7:0]  io_in_0_bits_req_inst,
  input  [63:0] io_in_0_bits_req_data,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_req_addr,
  input  [7:0]  io_in_1_bits_req_inst,
  input  [63:0] io_in_1_bits_req_data,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_req_addr,
  input  [7:0]  io_in_2_bits_req_inst,
  input  [63:0] io_in_2_bits_req_data,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_req_addr,
  input  [7:0]  io_in_3_bits_req_inst,
  input  [63:0] io_in_3_bits_req_data,
  output        io_in_4_ready,
  input         io_in_4_valid,
  input  [31:0] io_in_4_bits_req_addr,
  input  [7:0]  io_in_4_bits_req_inst,
  input  [63:0] io_in_4_bits_req_data,
  output        io_in_5_ready,
  input         io_in_5_valid,
  input  [31:0] io_in_5_bits_req_addr,
  input  [7:0]  io_in_5_bits_req_inst,
  input  [63:0] io_in_5_bits_req_data,
  output        io_in_6_ready,
  input         io_in_6_valid,
  input  [31:0] io_in_6_bits_req_addr,
  input  [7:0]  io_in_6_bits_req_inst,
  input  [63:0] io_in_6_bits_req_data,
  output        io_in_7_ready,
  input         io_in_7_valid,
  input  [31:0] io_in_7_bits_req_addr,
  input  [7:0]  io_in_7_bits_req_inst,
  input  [63:0] io_in_7_bits_req_data,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [7:0]  io_out_bits_req_inst,
  output [63:0] io_out_bits_req_data,
  output [2:0]  io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_7 = 3'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  wire [31:0] _GEN_9 = 3'h1 == io_chosen ? io_in_1_bits_req_addr : io_in_0_bits_req_addr; // @[Arbiter.scala 41:16]
  wire [7:0] _GEN_10 = 3'h1 == io_chosen ? io_in_1_bits_req_inst : io_in_0_bits_req_inst; // @[Arbiter.scala 41:16]
  wire [63:0] _GEN_11 = 3'h1 == io_chosen ? io_in_1_bits_req_data : io_in_0_bits_req_data; // @[Arbiter.scala 41:16]
  wire  _GEN_13 = 3'h2 == io_chosen ? io_in_2_valid : _GEN_7; // @[Arbiter.scala 41:16]
  wire [31:0] _GEN_15 = 3'h2 == io_chosen ? io_in_2_bits_req_addr : _GEN_9; // @[Arbiter.scala 41:16]
  wire [7:0] _GEN_16 = 3'h2 == io_chosen ? io_in_2_bits_req_inst : _GEN_10; // @[Arbiter.scala 41:16]
  wire [63:0] _GEN_17 = 3'h2 == io_chosen ? io_in_2_bits_req_data : _GEN_11; // @[Arbiter.scala 41:16]
  wire  _GEN_19 = 3'h3 == io_chosen ? io_in_3_valid : _GEN_13; // @[Arbiter.scala 41:16]
  wire [31:0] _GEN_21 = 3'h3 == io_chosen ? io_in_3_bits_req_addr : _GEN_15; // @[Arbiter.scala 41:16]
  wire [7:0] _GEN_22 = 3'h3 == io_chosen ? io_in_3_bits_req_inst : _GEN_16; // @[Arbiter.scala 41:16]
  wire [63:0] _GEN_23 = 3'h3 == io_chosen ? io_in_3_bits_req_data : _GEN_17; // @[Arbiter.scala 41:16]
  wire  _GEN_25 = 3'h4 == io_chosen ? io_in_4_valid : _GEN_19; // @[Arbiter.scala 41:16]
  wire [31:0] _GEN_27 = 3'h4 == io_chosen ? io_in_4_bits_req_addr : _GEN_21; // @[Arbiter.scala 41:16]
  wire [7:0] _GEN_28 = 3'h4 == io_chosen ? io_in_4_bits_req_inst : _GEN_22; // @[Arbiter.scala 41:16]
  wire [63:0] _GEN_29 = 3'h4 == io_chosen ? io_in_4_bits_req_data : _GEN_23; // @[Arbiter.scala 41:16]
  wire  _GEN_31 = 3'h5 == io_chosen ? io_in_5_valid : _GEN_25; // @[Arbiter.scala 41:16]
  wire [31:0] _GEN_33 = 3'h5 == io_chosen ? io_in_5_bits_req_addr : _GEN_27; // @[Arbiter.scala 41:16]
  wire [7:0] _GEN_34 = 3'h5 == io_chosen ? io_in_5_bits_req_inst : _GEN_28; // @[Arbiter.scala 41:16]
  wire [63:0] _GEN_35 = 3'h5 == io_chosen ? io_in_5_bits_req_data : _GEN_29; // @[Arbiter.scala 41:16]
  wire  _GEN_37 = 3'h6 == io_chosen ? io_in_6_valid : _GEN_31; // @[Arbiter.scala 41:16]
  wire [31:0] _GEN_39 = 3'h6 == io_chosen ? io_in_6_bits_req_addr : _GEN_33; // @[Arbiter.scala 41:16]
  wire [7:0] _GEN_40 = 3'h6 == io_chosen ? io_in_6_bits_req_inst : _GEN_34; // @[Arbiter.scala 41:16]
  wire [63:0] _GEN_41 = 3'h6 == io_chosen ? io_in_6_bits_req_data : _GEN_35; // @[Arbiter.scala 41:16]
  reg [2:0] lastGrant; // @[Reg.scala 15:16]
  wire  grantMask_1 = 3'h1 > lastGrant; // @[Arbiter.scala 67:49]
  wire  grantMask_2 = 3'h2 > lastGrant; // @[Arbiter.scala 67:49]
  wire  grantMask_3 = 3'h3 > lastGrant; // @[Arbiter.scala 67:49]
  wire  grantMask_4 = 3'h4 > lastGrant; // @[Arbiter.scala 67:49]
  wire  grantMask_5 = 3'h5 > lastGrant; // @[Arbiter.scala 67:49]
  wire  grantMask_6 = 3'h6 > lastGrant; // @[Arbiter.scala 67:49]
  wire  grantMask_7 = 3'h7 > lastGrant; // @[Arbiter.scala 67:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbiter.scala 68:75]
  wire  validMask_2 = io_in_2_valid & grantMask_2; // @[Arbiter.scala 68:75]
  wire  validMask_3 = io_in_3_valid & grantMask_3; // @[Arbiter.scala 68:75]
  wire  validMask_4 = io_in_4_valid & grantMask_4; // @[Arbiter.scala 68:75]
  wire  validMask_5 = io_in_5_valid & grantMask_5; // @[Arbiter.scala 68:75]
  wire  validMask_6 = io_in_6_valid & grantMask_6; // @[Arbiter.scala 68:75]
  wire  validMask_7 = io_in_7_valid & grantMask_7; // @[Arbiter.scala 68:75]
  wire  _T_2 = validMask_1 | validMask_2; // @[Arbiter.scala 31:68]
  wire  _T_3 = _T_2 | validMask_3; // @[Arbiter.scala 31:68]
  wire  _T_4 = _T_3 | validMask_4; // @[Arbiter.scala 31:68]
  wire  _T_5 = _T_4 | validMask_5; // @[Arbiter.scala 31:68]
  wire  _T_6 = _T_5 | validMask_6; // @[Arbiter.scala 31:68]
  wire  _T_7 = _T_6 | validMask_7; // @[Arbiter.scala 31:68]
  wire  _T_8 = _T_7 | io_in_0_valid; // @[Arbiter.scala 31:68]
  wire  _T_9 = _T_8 | io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  _T_10 = _T_9 | io_in_2_valid; // @[Arbiter.scala 31:68]
  wire  _T_11 = _T_10 | io_in_3_valid; // @[Arbiter.scala 31:68]
  wire  _T_12 = _T_11 | io_in_4_valid; // @[Arbiter.scala 31:68]
  wire  _T_13 = _T_12 | io_in_5_valid; // @[Arbiter.scala 31:68]
  wire  _T_14 = _T_13 | io_in_6_valid; // @[Arbiter.scala 31:68]
  wire  _T_16 = ~validMask_1; // @[Arbiter.scala 31:78]
  wire  _T_17 = ~_T_2; // @[Arbiter.scala 31:78]
  wire  _T_18 = ~_T_3; // @[Arbiter.scala 31:78]
  wire  _T_19 = ~_T_4; // @[Arbiter.scala 31:78]
  wire  _T_20 = ~_T_5; // @[Arbiter.scala 31:78]
  wire  _T_21 = ~_T_6; // @[Arbiter.scala 31:78]
  wire  _T_23 = ~_T_8; // @[Arbiter.scala 31:78]
  wire  _T_24 = ~_T_9; // @[Arbiter.scala 31:78]
  wire  _T_25 = ~_T_10; // @[Arbiter.scala 31:78]
  wire  _T_26 = ~_T_11; // @[Arbiter.scala 31:78]
  wire  _T_27 = ~_T_12; // @[Arbiter.scala 31:78]
  wire  _T_28 = ~_T_13; // @[Arbiter.scala 31:78]
  wire  _T_29 = ~_T_14; // @[Arbiter.scala 31:78]
  wire  _T_34 = _T_16 & grantMask_2; // @[Arbiter.scala 72:34]
  wire  _T_36 = _T_17 & grantMask_3; // @[Arbiter.scala 72:34]
  wire  _T_38 = _T_18 & grantMask_4; // @[Arbiter.scala 72:34]
  wire  _T_40 = _T_19 & grantMask_5; // @[Arbiter.scala 72:34]
  wire  _T_42 = _T_20 & grantMask_6; // @[Arbiter.scala 72:34]
  wire  _T_44 = _T_21 & grantMask_7; // @[Arbiter.scala 72:34]
  wire [2:0] _GEN_49 = io_in_6_valid ? 3'h6 : 3'h7; // @[Arbiter.scala 77:27]
  wire [2:0] _GEN_50 = io_in_5_valid ? 3'h5 : _GEN_49; // @[Arbiter.scala 77:27]
  wire [2:0] _GEN_51 = io_in_4_valid ? 3'h4 : _GEN_50; // @[Arbiter.scala 77:27]
  wire [2:0] _GEN_52 = io_in_3_valid ? 3'h3 : _GEN_51; // @[Arbiter.scala 77:27]
  wire [2:0] _GEN_53 = io_in_2_valid ? 3'h2 : _GEN_52; // @[Arbiter.scala 77:27]
  wire [2:0] _GEN_54 = io_in_1_valid ? 3'h1 : _GEN_53; // @[Arbiter.scala 77:27]
  wire [2:0] _GEN_55 = io_in_0_valid ? 3'h0 : _GEN_54; // @[Arbiter.scala 77:27]
  wire [2:0] _GEN_56 = validMask_7 ? 3'h7 : _GEN_55; // @[Arbiter.scala 79:25]
  wire [2:0] _GEN_57 = validMask_6 ? 3'h6 : _GEN_56; // @[Arbiter.scala 79:25]
  wire [2:0] _GEN_58 = validMask_5 ? 3'h5 : _GEN_57; // @[Arbiter.scala 79:25]
  wire [2:0] _GEN_59 = validMask_4 ? 3'h4 : _GEN_58; // @[Arbiter.scala 79:25]
  wire [2:0] _GEN_60 = validMask_3 ? 3'h3 : _GEN_59; // @[Arbiter.scala 79:25]
  wire [2:0] _GEN_61 = validMask_2 ? 3'h2 : _GEN_60; // @[Arbiter.scala 79:25]
  assign io_in_0_ready = ~_T_7; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = grantMask_1 | _T_23; // @[Arbiter.scala 60:16]
  assign io_in_2_ready = _T_34 | _T_24; // @[Arbiter.scala 60:16]
  assign io_in_3_ready = _T_36 | _T_25; // @[Arbiter.scala 60:16]
  assign io_in_4_ready = _T_38 | _T_26; // @[Arbiter.scala 60:16]
  assign io_in_5_ready = _T_40 | _T_27; // @[Arbiter.scala 60:16]
  assign io_in_6_ready = _T_42 | _T_28; // @[Arbiter.scala 60:16]
  assign io_in_7_ready = _T_44 | _T_29; // @[Arbiter.scala 60:16]
  assign io_out_valid = 3'h7 == io_chosen ? io_in_7_valid : _GEN_37; // @[Arbiter.scala 41:16]
  assign io_out_bits_req_addr = 3'h7 == io_chosen ? io_in_7_bits_req_addr : _GEN_39; // @[Arbiter.scala 42:15]
  assign io_out_bits_req_inst = 3'h7 == io_chosen ? io_in_7_bits_req_inst : _GEN_40; // @[Arbiter.scala 42:15]
  assign io_out_bits_req_data = 3'h7 == io_chosen ? io_in_7_bits_req_data : _GEN_41; // @[Arbiter.scala 42:15]
  assign io_chosen = validMask_1 ? 3'h1 : _GEN_61; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_out_valid) begin
      lastGrant <= io_chosen;
    end
  end
endmodule
module Arbiter_4(
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_addr,
  input         io_in_4_valid,
  input  [31:0] io_in_4_bits_addr,
  input         io_in_5_valid,
  input  [31:0] io_in_5_bits_addr,
  input         io_in_6_valid,
  input  [31:0] io_in_6_bits_addr,
  input         io_in_7_valid,
  input  [31:0] io_in_7_bits_addr,
  input         io_in_8_valid,
  input  [31:0] io_in_8_bits_addr,
  output        io_out_valid,
  output [31:0] io_out_bits_addr
);
  wire [31:0] _GEN_2 = io_in_7_valid ? io_in_7_bits_addr : io_in_8_bits_addr; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_6 = io_in_6_valid ? io_in_6_bits_addr : _GEN_2; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_10 = io_in_5_valid ? io_in_5_bits_addr : _GEN_6; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_14 = io_in_4_valid ? io_in_4_bits_addr : _GEN_10; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_18 = io_in_3_valid ? io_in_3_bits_addr : _GEN_14; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_22 = io_in_2_valid ? io_in_2_bits_addr : _GEN_18; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_26 = io_in_1_valid ? io_in_1_bits_addr : _GEN_22; // @[Arbiter.scala 126:27]
  wire  _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  _T_1 = _T | io_in_2_valid; // @[Arbiter.scala 31:68]
  wire  _T_2 = _T_1 | io_in_3_valid; // @[Arbiter.scala 31:68]
  wire  _T_3 = _T_2 | io_in_4_valid; // @[Arbiter.scala 31:68]
  wire  _T_4 = _T_3 | io_in_5_valid; // @[Arbiter.scala 31:68]
  wire  _T_5 = _T_4 | io_in_6_valid; // @[Arbiter.scala 31:68]
  wire  _T_6 = _T_5 | io_in_7_valid; // @[Arbiter.scala 31:68]
  wire  grant_8 = ~_T_6; // @[Arbiter.scala 31:78]
  wire  _T_16 = ~grant_8; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_16 | io_in_8_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_26; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
endmodule
module Arbiter_5(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [1:0]  io_in_0_bits_event,
  input  [31:0] io_in_0_bits_addr,
  input  [63:0] io_in_0_bits_data,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [1:0]  io_in_1_bits_event,
  input  [31:0] io_in_1_bits_addr,
  input  [63:0] io_in_1_bits_data,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [1:0]  io_in_2_bits_event,
  input  [31:0] io_in_2_bits_addr,
  input  [63:0] io_in_2_bits_data,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [1:0]  io_in_3_bits_event,
  input  [31:0] io_in_3_bits_addr,
  input  [63:0] io_in_3_bits_data,
  output        io_in_4_ready,
  input         io_in_4_valid,
  input  [1:0]  io_in_4_bits_event,
  input  [31:0] io_in_4_bits_addr,
  input  [63:0] io_in_4_bits_data,
  output        io_in_5_ready,
  input         io_in_5_valid,
  input  [1:0]  io_in_5_bits_event,
  input  [31:0] io_in_5_bits_addr,
  input  [63:0] io_in_5_bits_data,
  output        io_in_6_ready,
  input         io_in_6_valid,
  input  [1:0]  io_in_6_bits_event,
  input  [31:0] io_in_6_bits_addr,
  input  [63:0] io_in_6_bits_data,
  output        io_in_7_ready,
  input         io_in_7_valid,
  input  [1:0]  io_in_7_bits_event,
  input  [31:0] io_in_7_bits_addr,
  input  [63:0] io_in_7_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output [1:0]  io_out_bits_event,
  output [31:0] io_out_bits_addr,
  output [63:0] io_out_bits_data
);
  wire [63:0] _GEN_1 = io_in_6_valid ? io_in_6_bits_data : io_in_7_bits_data; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_2 = io_in_6_valid ? io_in_6_bits_addr : io_in_7_bits_addr; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_3 = io_in_6_valid ? io_in_6_bits_event : io_in_7_bits_event; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_5 = io_in_5_valid ? io_in_5_bits_data : _GEN_1; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_6 = io_in_5_valid ? io_in_5_bits_addr : _GEN_2; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_7 = io_in_5_valid ? io_in_5_bits_event : _GEN_3; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_9 = io_in_4_valid ? io_in_4_bits_data : _GEN_5; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_10 = io_in_4_valid ? io_in_4_bits_addr : _GEN_6; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_11 = io_in_4_valid ? io_in_4_bits_event : _GEN_7; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_13 = io_in_3_valid ? io_in_3_bits_data : _GEN_9; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_14 = io_in_3_valid ? io_in_3_bits_addr : _GEN_10; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_15 = io_in_3_valid ? io_in_3_bits_event : _GEN_11; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_17 = io_in_2_valid ? io_in_2_bits_data : _GEN_13; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_18 = io_in_2_valid ? io_in_2_bits_addr : _GEN_14; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_19 = io_in_2_valid ? io_in_2_bits_event : _GEN_15; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_21 = io_in_1_valid ? io_in_1_bits_data : _GEN_17; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_22 = io_in_1_valid ? io_in_1_bits_addr : _GEN_18; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_23 = io_in_1_valid ? io_in_1_bits_event : _GEN_19; // @[Arbiter.scala 126:27]
  wire  _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  _T_1 = _T | io_in_2_valid; // @[Arbiter.scala 31:68]
  wire  _T_2 = _T_1 | io_in_3_valid; // @[Arbiter.scala 31:68]
  wire  _T_3 = _T_2 | io_in_4_valid; // @[Arbiter.scala 31:68]
  wire  _T_4 = _T_3 | io_in_5_valid; // @[Arbiter.scala 31:68]
  wire  _T_5 = _T_4 | io_in_6_valid; // @[Arbiter.scala 31:68]
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  grant_2 = ~_T; // @[Arbiter.scala 31:78]
  wire  grant_3 = ~_T_1; // @[Arbiter.scala 31:78]
  wire  grant_4 = ~_T_2; // @[Arbiter.scala 31:78]
  wire  grant_5 = ~_T_3; // @[Arbiter.scala 31:78]
  wire  grant_6 = ~_T_4; // @[Arbiter.scala 31:78]
  wire  grant_7 = ~_T_5; // @[Arbiter.scala 31:78]
  wire  _T_14 = ~grant_7; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_2_ready = grant_2 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_3_ready = grant_3 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_4_ready = grant_4 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_5_ready = grant_5 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_6_ready = grant_6 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_7_ready = grant_7 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_14 | io_in_7_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_event = io_in_0_valid ? io_in_0_bits_event : _GEN_23; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_22; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : _GEN_21; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
endmodule
module Queue_7(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_inst_event,
  input  [31:0] io_enq_bits_inst_addr,
  input  [63:0] io_enq_bits_inst_data,
  input  [1:0]  io_enq_bits_tbeOut_state_state,
  input  [2:0]  io_enq_bits_tbeOut_way,
  input  [31:0] io_enq_bits_tbeOut_fields_0,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_inst_event,
  output [31:0] io_deq_bits_inst_addr,
  output [63:0] io_deq_bits_inst_data,
  output [1:0]  io_deq_bits_tbeOut_state_state,
  output [2:0]  io_deq_bits_tbeOut_way,
  output [31:0] io_deq_bits_tbeOut_fields_0
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_inst_event [0:0]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_inst_event__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_inst_event__T_7_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_inst_event__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst_event__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst_event__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst_event__T_3_en; // @[Decoupled.scala 209:16]
  reg [31:0] ram_inst_addr [0:0]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_inst_addr__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_inst_addr__T_7_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_inst_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_inst_data [0:0]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_inst_data__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_inst_data__T_7_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_inst_data__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [1:0] ram_tbeOut_state_state [0:0]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_tbeOut_state_state__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_state_state__T_7_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_tbeOut_state_state__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_state_state__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_state_state__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_state_state__T_3_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_tbeOut_way [0:0]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_tbeOut_way__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_way__T_7_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_tbeOut_way__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_way__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_way__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_way__T_3_en; // @[Decoupled.scala 209:16]
  reg [31:0] ram_tbeOut_fields_0 [0:0]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_tbeOut_fields_0__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_fields_0__T_7_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_tbeOut_fields_0__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_fields_0__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_fields_0__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_fields_0__T_3_en; // @[Decoupled.scala 209:16]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram_inst_event__T_7_addr = 1'h0;
  assign ram_inst_event__T_7_data = ram_inst_event[ram_inst_event__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst_event__T_3_data = io_enq_bits_inst_event;
  assign ram_inst_event__T_3_addr = 1'h0;
  assign ram_inst_event__T_3_mask = 1'h1;
  assign ram_inst_event__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst_addr__T_7_addr = 1'h0;
  assign ram_inst_addr__T_7_data = ram_inst_addr[ram_inst_addr__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst_addr__T_3_data = io_enq_bits_inst_addr;
  assign ram_inst_addr__T_3_addr = 1'h0;
  assign ram_inst_addr__T_3_mask = 1'h1;
  assign ram_inst_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst_data__T_7_addr = 1'h0;
  assign ram_inst_data__T_7_data = ram_inst_data[ram_inst_data__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst_data__T_3_data = io_enq_bits_inst_data;
  assign ram_inst_data__T_3_addr = 1'h0;
  assign ram_inst_data__T_3_mask = 1'h1;
  assign ram_inst_data__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_tbeOut_state_state__T_7_addr = 1'h0;
  assign ram_tbeOut_state_state__T_7_data = ram_tbeOut_state_state[ram_tbeOut_state_state__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_tbeOut_state_state__T_3_data = io_enq_bits_tbeOut_state_state;
  assign ram_tbeOut_state_state__T_3_addr = 1'h0;
  assign ram_tbeOut_state_state__T_3_mask = 1'h1;
  assign ram_tbeOut_state_state__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_tbeOut_way__T_7_addr = 1'h0;
  assign ram_tbeOut_way__T_7_data = ram_tbeOut_way[ram_tbeOut_way__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_tbeOut_way__T_3_data = io_enq_bits_tbeOut_way;
  assign ram_tbeOut_way__T_3_addr = 1'h0;
  assign ram_tbeOut_way__T_3_mask = 1'h1;
  assign ram_tbeOut_way__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_tbeOut_fields_0__T_7_addr = 1'h0;
  assign ram_tbeOut_fields_0__T_7_data = ram_tbeOut_fields_0[ram_tbeOut_fields_0__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_tbeOut_fields_0__T_3_data = io_enq_bits_tbeOut_fields_0;
  assign ram_tbeOut_fields_0__T_3_addr = 1'h0;
  assign ram_tbeOut_fields_0__T_3_mask = 1'h1;
  assign ram_tbeOut_fields_0__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_inst_event = ram_inst_event__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst_addr = ram_inst_addr__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst_data = ram_inst_data__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_tbeOut_state_state = ram_tbeOut_state_state__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_tbeOut_way = ram_tbeOut_way__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_tbeOut_fields_0 = ram_tbeOut_fields_0__T_7_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_inst_event[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_inst_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_inst_data[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tbeOut_state_state[initvar] = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tbeOut_way[initvar] = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tbeOut_fields_0[initvar] = _RAND_5[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  maybe_full = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_inst_event__T_3_en & ram_inst_event__T_3_mask) begin
      ram_inst_event[ram_inst_event__T_3_addr] <= ram_inst_event__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst_addr__T_3_en & ram_inst_addr__T_3_mask) begin
      ram_inst_addr[ram_inst_addr__T_3_addr] <= ram_inst_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst_data__T_3_en & ram_inst_data__T_3_mask) begin
      ram_inst_data[ram_inst_data__T_3_addr] <= ram_inst_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_tbeOut_state_state__T_3_en & ram_tbeOut_state_state__T_3_mask) begin
      ram_tbeOut_state_state[ram_tbeOut_state_state__T_3_addr] <= ram_tbeOut_state_state__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_tbeOut_way__T_3_en & ram_tbeOut_way__T_3_mask) begin
      ram_tbeOut_way[ram_tbeOut_way__T_3_addr] <= ram_tbeOut_way__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_tbeOut_fields_0__T_3_en & ram_tbeOut_fields_0__T_3_mask) begin
      ram_tbeOut_fields_0[ram_tbeOut_fields_0__T_3_addr] <= ram_tbeOut_fields_0__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_4) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_8(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_event,
  input  [31:0] io_enq_bits_addr,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_event,
  output [31:0] io_deq_bits_addr,
  output [63:0] io_deq_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_event [0:0]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_event__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_event__T_7_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_event__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_event__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_event__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_event__T_3_en; // @[Decoupled.scala 209:16]
  reg [31:0] ram_addr [0:0]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_7_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:0]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_7_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram_event__T_7_addr = 1'h0;
  assign ram_event__T_7_data = ram_event[ram_event__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_event__T_3_data = io_enq_bits_event;
  assign ram_event__T_3_addr = 1'h0;
  assign ram_event__T_3_mask = 1'h1;
  assign ram_event__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_addr__T_7_addr = 1'h0;
  assign ram_addr__T_7_data = ram_addr[ram_addr__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_3_data = io_enq_bits_addr;
  assign ram_addr__T_3_addr = 1'h0;
  assign ram_addr__T_3_mask = 1'h1;
  assign ram_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_7_addr = 1'h0;
  assign ram_data__T_7_data = ram_data[ram_data__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = 1'h0;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_event = ram_event__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_addr = ram_addr__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_7_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_event[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_event__T_3_en & ram_event__T_3_mask) begin
      ram_event[ram_event__T_3_addr] <= ram_event__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_addr__T_3_en & ram_addr__T_3_mask) begin
      ram_addr[ram_addr__T_3_addr] <= ram_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_4) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_17(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_inst,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_inst,
  output [63:0] io_deq_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:0]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_7_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [7:0] ram_inst [0:0]; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_7_addr; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:0]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_7_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram_addr__T_7_addr = 1'h0;
  assign ram_addr__T_7_data = ram_addr[ram_addr__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_3_data = io_enq_bits_addr;
  assign ram_addr__T_3_addr = 1'h0;
  assign ram_addr__T_3_mask = 1'h1;
  assign ram_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst__T_7_addr = 1'h0;
  assign ram_inst__T_7_data = ram_inst[ram_inst__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst__T_3_data = io_enq_bits_inst;
  assign ram_inst__T_3_addr = 1'h0;
  assign ram_inst__T_3_mask = 1'h1;
  assign ram_inst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_7_addr = 1'h0;
  assign ram_data__T_7_data = ram_data[ram_data__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = 1'h0;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst = ram_inst__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_7_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_inst[initvar] = _RAND_1[7:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_3_en & ram_addr__T_3_mask) begin
      ram_addr[ram_addr__T_3_addr] <= ram_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst__T_3_en & ram_inst__T_3_mask) begin
      ram_inst[ram_inst__T_3_addr] <= ram_inst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_4) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_33(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [1:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [1:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram [0:0]; // @[Decoupled.scala 209:16]
  wire [1:0] ram__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram__T_7_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram__T_3_en; // @[Decoupled.scala 209:16]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  _T_1 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = io_deq_ready ? 1'h0 : _T_1; // @[Decoupled.scala 240:27]
  wire  do_enq = empty ? _GEN_7 : _T_1; // @[Decoupled.scala 237:18]
  wire  do_deq = empty ? 1'h0 : _T_2; // @[Decoupled.scala 237:18]
  wire  _T_4 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  wire  _T_5 = ~empty; // @[Decoupled.scala 231:19]
  assign ram__T_7_addr = 1'h0;
  assign ram__T_7_data = ram[ram__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram__T_3_data = io_enq_bits;
  assign ram__T_3_addr = 1'h0;
  assign ram__T_3_mask = 1'h1;
  assign ram__T_3_en = empty ? _GEN_7 : _T_1;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = io_enq_valid | _T_5; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits = empty ? io_enq_bits : ram__T_7_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maybe_full = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_3_en & ram__T_3_mask) begin
      ram[ram__T_3_addr] <= ram__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_4) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _T_1;
        end
      end else begin
        maybe_full <= _T_1;
      end
    end
  end
endmodule
module Queue_35(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] ram [0:0]; // @[Decoupled.scala 209:16]
  wire [15:0] ram__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram__T_7_addr; // @[Decoupled.scala 209:16]
  wire [15:0] ram__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram__T_3_en; // @[Decoupled.scala 209:16]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram__T_7_addr = 1'h0;
  assign ram__T_7_data = ram[ram__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram__T_3_data = io_enq_bits;
  assign ram__T_3_addr = 1'h0;
  assign ram__T_3_mask = 1'h1;
  assign ram__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits = ram__T_7_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maybe_full = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_3_en & ram__T_3_mask) begin
      ram[ram__T_3_addr] <= ram__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_4) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_36(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [1:0]  io_enq_bits_way,
  input  [63:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_replaceWay,
  input  [31:0] io_enq_bits_tbeFields_0,
  input  [27:0] io_enq_bits_action_signals,
  input  [3:0]  io_enq_bits_action_actionType,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [1:0]  io_deq_bits_way,
  output [63:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_replaceWay,
  output [31:0] io_deq_bits_tbeFields_0,
  output [27:0] io_deq_bits_action_signals,
  output [3:0]  io_deq_bits_action_actionType
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:0]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_33_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_27_en; // @[Decoupled.scala 209:16]
  reg [1:0] ram_way [0:0]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_way__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_way__T_33_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_way__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_way__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_way__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_way__T_27_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:0]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_33_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_27_en; // @[Decoupled.scala 209:16]
  reg [1:0] ram_replaceWay [0:0]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_replaceWay__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_replaceWay__T_33_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_replaceWay__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_replaceWay__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_replaceWay__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_replaceWay__T_27_en; // @[Decoupled.scala 209:16]
  reg [31:0] ram_tbeFields_0 [0:0]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_tbeFields_0__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeFields_0__T_33_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_tbeFields_0__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeFields_0__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_tbeFields_0__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_tbeFields_0__T_27_en; // @[Decoupled.scala 209:16]
  reg [27:0] ram_action_signals [0:0]; // @[Decoupled.scala 209:16]
  wire [27:0] ram_action_signals__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_action_signals__T_33_addr; // @[Decoupled.scala 209:16]
  wire [27:0] ram_action_signals__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_action_signals__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_action_signals__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_action_signals__T_27_en; // @[Decoupled.scala 209:16]
  reg [3:0] ram_action_actionType [0:0]; // @[Decoupled.scala 209:16]
  wire [3:0] ram_action_actionType__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_action_actionType__T_33_addr; // @[Decoupled.scala 209:16]
  wire [3:0] ram_action_actionType__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_action_actionType__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_action_actionType__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_action_actionType__T_27_en; // @[Decoupled.scala 209:16]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = do_enq != io_deq_valid; // @[Decoupled.scala 227:16]
  assign ram_addr__T_33_addr = 1'h0;
  assign ram_addr__T_33_data = ram_addr[ram_addr__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_27_data = io_enq_bits_addr;
  assign ram_addr__T_27_addr = 1'h0;
  assign ram_addr__T_27_mask = 1'h1;
  assign ram_addr__T_27_en = io_enq_ready & io_enq_valid;
  assign ram_way__T_33_addr = 1'h0;
  assign ram_way__T_33_data = ram_way[ram_way__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_way__T_27_data = io_enq_bits_way;
  assign ram_way__T_27_addr = 1'h0;
  assign ram_way__T_27_mask = 1'h1;
  assign ram_way__T_27_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_33_addr = 1'h0;
  assign ram_data__T_33_data = ram_data[ram_data__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_27_data = io_enq_bits_data;
  assign ram_data__T_27_addr = 1'h0;
  assign ram_data__T_27_mask = 1'h1;
  assign ram_data__T_27_en = io_enq_ready & io_enq_valid;
  assign ram_replaceWay__T_33_addr = 1'h0;
  assign ram_replaceWay__T_33_data = ram_replaceWay[ram_replaceWay__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_replaceWay__T_27_data = io_enq_bits_replaceWay;
  assign ram_replaceWay__T_27_addr = 1'h0;
  assign ram_replaceWay__T_27_mask = 1'h1;
  assign ram_replaceWay__T_27_en = io_enq_ready & io_enq_valid;
  assign ram_tbeFields_0__T_33_addr = 1'h0;
  assign ram_tbeFields_0__T_33_data = ram_tbeFields_0[ram_tbeFields_0__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_tbeFields_0__T_27_data = io_enq_bits_tbeFields_0;
  assign ram_tbeFields_0__T_27_addr = 1'h0;
  assign ram_tbeFields_0__T_27_mask = 1'h1;
  assign ram_tbeFields_0__T_27_en = io_enq_ready & io_enq_valid;
  assign ram_action_signals__T_33_addr = 1'h0;
  assign ram_action_signals__T_33_data = ram_action_signals[ram_action_signals__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_action_signals__T_27_data = io_enq_bits_action_signals;
  assign ram_action_signals__T_27_addr = 1'h0;
  assign ram_action_signals__T_27_mask = 1'h1;
  assign ram_action_signals__T_27_en = io_enq_ready & io_enq_valid;
  assign ram_action_actionType__T_33_addr = 1'h0;
  assign ram_action_actionType__T_33_data = ram_action_actionType[ram_action_actionType__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_action_actionType__T_27_data = io_enq_bits_action_actionType;
  assign ram_action_actionType__T_27_addr = 1'h0;
  assign ram_action_actionType__T_27_mask = 1'h1;
  assign ram_action_actionType__T_27_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = 1'h1; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_33_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_way = ram_way__T_33_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_33_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_replaceWay = ram_replaceWay__T_33_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_tbeFields_0 = ram_tbeFields_0__T_33_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_action_signals = ram_action_signals__T_33_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_action_actionType = ram_action_actionType__T_33_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_way[initvar] = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_replaceWay[initvar] = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tbeFields_0[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_action_signals[initvar] = _RAND_5[27:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_action_actionType[initvar] = _RAND_6[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_27_en & ram_addr__T_27_mask) begin
      ram_addr[ram_addr__T_27_addr] <= ram_addr__T_27_data; // @[Decoupled.scala 209:16]
    end
    if(ram_way__T_27_en & ram_way__T_27_mask) begin
      ram_way[ram_way__T_27_addr] <= ram_way__T_27_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_27_en & ram_data__T_27_mask) begin
      ram_data[ram_data__T_27_addr] <= ram_data__T_27_data; // @[Decoupled.scala 209:16]
    end
    if(ram_replaceWay__T_27_en & ram_replaceWay__T_27_mask) begin
      ram_replaceWay[ram_replaceWay__T_27_addr] <= ram_replaceWay__T_27_data; // @[Decoupled.scala 209:16]
    end
    if(ram_tbeFields_0__T_27_en & ram_tbeFields_0__T_27_mask) begin
      ram_tbeFields_0[ram_tbeFields_0__T_27_addr] <= ram_tbeFields_0__T_27_data; // @[Decoupled.scala 209:16]
    end
    if(ram_action_signals__T_27_en & ram_action_signals__T_27_mask) begin
      ram_action_signals[ram_action_signals__T_27_addr] <= ram_action_signals__T_27_data; // @[Decoupled.scala 209:16]
    end
    if(ram_action_actionType__T_27_en & ram_action_actionType__T_27_mask) begin
      ram_action_actionType[ram_action_actionType__T_27_addr] <= ram_action_actionType__T_27_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_30) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module MIMOQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_0_way,
  input  [31:0] io_enq_bits_0_addr,
  input  [1:0]  io_enq_bits_1_way,
  input  [31:0] io_enq_bits_1_addr,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_0_way,
  output [31:0] io_deq_bits_0_addr,
  output [3:0]  io_count
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_way [0:7]; // @[MIMOQueue.scala 56:16]
  wire [1:0] ram_way__T_22_data; // @[MIMOQueue.scala 56:16]
  wire [2:0] ram_way__T_22_addr; // @[MIMOQueue.scala 56:16]
  wire [1:0] ram_way__T_7_data; // @[MIMOQueue.scala 56:16]
  wire [2:0] ram_way__T_7_addr; // @[MIMOQueue.scala 56:16]
  wire  ram_way__T_7_mask; // @[MIMOQueue.scala 56:16]
  wire  ram_way__T_7_en; // @[MIMOQueue.scala 56:16]
  wire [1:0] ram_way__T_10_data; // @[MIMOQueue.scala 56:16]
  wire [2:0] ram_way__T_10_addr; // @[MIMOQueue.scala 56:16]
  wire  ram_way__T_10_mask; // @[MIMOQueue.scala 56:16]
  wire  ram_way__T_10_en; // @[MIMOQueue.scala 56:16]
  reg [31:0] ram_addr [0:7]; // @[MIMOQueue.scala 56:16]
  wire [31:0] ram_addr__T_22_data; // @[MIMOQueue.scala 56:16]
  wire [2:0] ram_addr__T_22_addr; // @[MIMOQueue.scala 56:16]
  wire [31:0] ram_addr__T_7_data; // @[MIMOQueue.scala 56:16]
  wire [2:0] ram_addr__T_7_addr; // @[MIMOQueue.scala 56:16]
  wire  ram_addr__T_7_mask; // @[MIMOQueue.scala 56:16]
  wire  ram_addr__T_7_en; // @[MIMOQueue.scala 56:16]
  wire [31:0] ram_addr__T_10_data; // @[MIMOQueue.scala 56:16]
  wire [2:0] ram_addr__T_10_addr; // @[MIMOQueue.scala 56:16]
  wire  ram_addr__T_10_mask; // @[MIMOQueue.scala 56:16]
  wire  ram_addr__T_10_en; // @[MIMOQueue.scala 56:16]
  reg [2:0] value; // @[Counter.scala 29:33]
  reg [2:0] value_1; // @[Counter.scala 29:33]
  reg  maybe_full; // @[MIMOQueue.scala 59:27]
  wire  ptr_match = value == value_1; // @[MIMOQueue.scala 62:33]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _T_5 = {{1'd0}, value}; // @[MIMOQueue.scala 77:25]
  wire [2:0] _T_12 = value + 3'h2; // @[MIMOQueue.scala 79:36]
  wire [2:0] _T_14 = value_1 + 3'h1; // @[MIMOQueue.scala 86:36]
  wire  _T_15 = do_enq != io_deq_valid; // @[MIMOQueue.scala 91:16]
  wire [2:0] ptr_diff = value - value_1; // @[MIMOQueue.scala 97:32]
  wire  _T_18 = io_count > 4'h0; // @[MIMOQueue.scala 100:18]
  wire [3:0] _T_20 = {{1'd0}, value_1}; // @[MIMOQueue.scala 106:73]
  wire  _T_25 = maybe_full & ptr_match; // @[MIMOQueue.scala 123:32]
  assign ram_way__T_22_addr = _T_20[2:0];
  assign ram_way__T_22_data = ram_way[ram_way__T_22_addr]; // @[MIMOQueue.scala 56:16]
  assign ram_way__T_7_data = io_enq_bits_0_way;
  assign ram_way__T_7_addr = _T_5[2:0];
  assign ram_way__T_7_mask = 1'h1;
  assign ram_way__T_7_en = io_enq_ready & io_enq_valid;
  assign ram_way__T_10_data = io_enq_bits_1_way;
  assign ram_way__T_10_addr = value + 3'h1;
  assign ram_way__T_10_mask = 1'h1;
  assign ram_way__T_10_en = io_enq_ready & io_enq_valid;
  assign ram_addr__T_22_addr = _T_20[2:0];
  assign ram_addr__T_22_data = ram_addr[ram_addr__T_22_addr]; // @[MIMOQueue.scala 56:16]
  assign ram_addr__T_7_data = io_enq_bits_0_addr;
  assign ram_addr__T_7_addr = _T_5[2:0];
  assign ram_addr__T_7_mask = 1'h1;
  assign ram_addr__T_7_en = io_enq_ready & io_enq_valid;
  assign ram_addr__T_10_data = io_enq_bits_1_addr;
  assign ram_addr__T_10_addr = value + 3'h1;
  assign ram_addr__T_10_mask = 1'h1;
  assign ram_addr__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = 1'h1; // @[MIMOQueue.scala 95:16 MIMOQueue.scala 119:40]
  assign io_deq_valid = io_count > 4'h0; // @[MIMOQueue.scala 101:18 MIMOQueue.scala 103:18]
  assign io_deq_bits_0_way = _T_18 ? ram_way__T_22_data : 2'h0; // @[MIMOQueue.scala 106:20]
  assign io_deq_bits_0_addr = _T_18 ? ram_addr__T_22_data : 32'h0; // @[MIMOQueue.scala 106:20]
  assign io_count = _T_25 ? 4'h8 : {{1'd0}, ptr_diff}; // @[MIMOQueue.scala 123:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_way[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_way__T_7_en & ram_way__T_7_mask) begin
      ram_way[ram_way__T_7_addr] <= ram_way__T_7_data; // @[MIMOQueue.scala 56:16]
    end
    if(ram_way__T_10_en & ram_way__T_10_mask) begin
      ram_way[ram_way__T_10_addr] <= ram_way__T_10_data; // @[MIMOQueue.scala 56:16]
    end
    if(ram_addr__T_7_en & ram_addr__T_7_mask) begin
      ram_addr[ram_addr__T_7_addr] <= ram_addr__T_7_data; // @[MIMOQueue.scala 56:16]
    end
    if(ram_addr__T_10_en & ram_addr__T_10_mask) begin
      ram_addr[ram_addr__T_10_addr] <= ram_addr__T_10_data; // @[MIMOQueue.scala 56:16]
    end
    if (reset) begin
      value <= 3'h0;
    end else if (do_enq) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else if (io_deq_valid) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_15) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Computation(
  input         clock,
  input         reset,
  input         io_instruction_valid,
  input  [27:0] io_instruction_bits,
  input         io_clear,
  input         io_op1_valid,
  input  [63:0] io_op1_bits,
  input         io_op2_valid,
  input  [63:0] io_op2_bits,
  output [15:0] io_pc,
  output [63:0] io_reg_file_0,
  output [63:0] io_reg_file_1,
  output [63:0] io_reg_file_2,
  output [63:0] io_reg_file_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] function_ = io_instruction_bits[3:0]; // @[Computation.scala 69:42]
  wire [5:0] write_addr = io_instruction_bits[9:4]; // @[Computation.scala 70:42]
  wire [1:0] read_addr1 = io_instruction_bits[11:10]; // @[Computation.scala 73:42]
  wire [15:0] read_addr2 = io_instruction_bits[27:12]; // @[Computation.scala 74:42]
  reg [63:0] reg_file_3; // @[Computation.scala 86:27]
  reg [63:0] reg_file_2; // @[Computation.scala 86:27]
  reg [63:0] reg_file_1; // @[Computation.scala 86:27]
  reg [63:0] reg_file_0; // @[Computation.scala 86:27]
  wire [63:0] _GEN_13 = 2'h1 == read_addr1 ? reg_file_1 : reg_file_0; // @[Computation.scala 92:14]
  wire [63:0] _GEN_14 = 2'h2 == read_addr1 ? reg_file_2 : _GEN_13; // @[Computation.scala 92:14]
  wire [63:0] reg_out1 = 2'h3 == read_addr1 ? reg_file_3 : _GEN_14; // @[Computation.scala 92:14]
  wire [63:0] alu_in1 = io_op1_valid ? io_op1_bits : reg_out1; // @[Computation.scala 82:19]
  wire [63:0] _GEN_17 = 2'h1 == read_addr2[1:0] ? reg_file_1 : reg_file_0; // @[Computation.scala 93:14]
  wire [63:0] _GEN_18 = 2'h2 == read_addr2[1:0] ? reg_file_2 : _GEN_17; // @[Computation.scala 93:14]
  wire [63:0] reg_out2 = 2'h3 == read_addr2[1:0] ? reg_file_3 : _GEN_18; // @[Computation.scala 93:14]
  wire [63:0] alu_in2 = io_op2_valid ? io_op2_bits : reg_out2; // @[Computation.scala 83:19]
  wire  _T_3 = function_ != 4'h6; // @[Computation.scala 88:55]
  wire  _T_4 = function_ != 4'h7; // @[Computation.scala 88:75]
  wire  _T_5 = _T_3 & _T_4; // @[Computation.scala 88:63]
  wire  write_en = io_instruction_valid & _T_5; // @[Computation.scala 88:42]
  wire  _T_10 = 4'h0 == function_; // @[Conditional.scala 37:30]
  wire [63:0] _T_12 = alu_in1 + alu_in2; // @[Computation.scala 33:38]
  wire  _T_13 = 4'h1 == function_; // @[Conditional.scala 37:30]
  wire [63:0] _T_14 = alu_in1 & alu_in2; // @[Computation.scala 34:38]
  wire  _T_15 = 4'h2 == function_; // @[Conditional.scala 37:30]
  wire [63:0] _T_17 = alu_in1 - alu_in2; // @[Computation.scala 35:38]
  wire  _T_18 = 4'h3 == function_; // @[Conditional.scala 37:30]
  wire [63:0] _T_19 = alu_in1 >> alu_in2; // @[Computation.scala 36:42]
  wire  _T_20 = 4'h4 == function_; // @[Conditional.scala 37:30]
  wire [318:0] _GEN_29 = {{255'd0}, alu_in1}; // @[Computation.scala 37:42]
  wire [318:0] _T_22 = _GEN_29 << alu_in2[7:0]; // @[Computation.scala 37:42]
  wire  _T_23 = 4'h5 == function_; // @[Conditional.scala 37:30]
  wire [63:0] _T_24 = alu_in1 ^ alu_in2; // @[Computation.scala 38:38]
  wire  _T_25 = 4'h6 == function_; // @[Conditional.scala 37:30]
  wire  _T_26 = alu_in1 < alu_in2; // @[Computation.scala 39:43]
  wire [63:0] _T_8 = {{58'd0}, write_addr}; // @[Computation.scala 97:93 Computation.scala 97:93]
  wire [63:0] _T_27 = _T_26 ? _T_8 : 64'h0; // @[Computation.scala 39:38]
  wire  _T_28 = 4'h7 == function_; // @[Conditional.scala 37:30]
  wire  _T_29 = alu_in1 != alu_in2; // @[Computation.scala 40:43]
  wire [63:0] _T_30 = _T_29 ? _T_8 : 64'h0; // @[Computation.scala 40:38]
  wire  _T_31 = 4'h8 == function_; // @[Conditional.scala 37:30]
  wire [63:0] _T_32 = alu_in1 | alu_in2; // @[Computation.scala 41:37]
  wire [63:0] _GEN_20 = _T_31 ? _T_32 : 64'h0; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_21 = _T_28 ? _T_30 : _GEN_20; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_22 = _T_25 ? _T_27 : _GEN_21; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_23 = _T_23 ? _T_24 : _GEN_22; // @[Conditional.scala 39:67]
  wire [318:0] _GEN_24 = _T_20 ? _T_22 : {{255'd0}, _GEN_23}; // @[Conditional.scala 39:67]
  wire [318:0] _GEN_25 = _T_18 ? {{255'd0}, _T_19} : _GEN_24; // @[Conditional.scala 39:67]
  wire [318:0] _GEN_26 = _T_15 ? {{255'd0}, _T_17} : _GEN_25; // @[Conditional.scala 39:67]
  wire [318:0] _GEN_27 = _T_13 ? {{255'd0}, _T_14} : _GEN_26; // @[Conditional.scala 39:67]
  wire [318:0] _GEN_28 = _T_10 ? {{255'd0}, _T_12} : _GEN_27; // @[Conditional.scala 40:58]
  wire [63:0] result = io_instruction_valid ? _GEN_28[63:0] : 64'h0; // @[Computation.scala 97:18]
  assign io_pc = _T_5 ? 16'h0 : result[15:0]; // @[Computation.scala 98:11]
  assign io_reg_file_0 = reg_file_0; // @[Computation.scala 94:17]
  assign io_reg_file_1 = reg_file_1; // @[Computation.scala 94:17]
  assign io_reg_file_2 = reg_file_2; // @[Computation.scala 94:17]
  assign io_reg_file_3 = reg_file_3; // @[Computation.scala 94:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  reg_file_3 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  reg_file_2 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  reg_file_1 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  reg_file_0 = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      reg_file_3 <= 64'h0;
    end else if (io_clear) begin
      reg_file_3 <= 64'h0;
    end else if (write_en) begin
      if (2'h3 == write_addr[1:0]) begin
        if (io_instruction_valid) begin
          reg_file_3 <= _GEN_28[63:0];
        end else begin
          reg_file_3 <= 64'h0;
        end
      end
    end
    if (reset) begin
      reg_file_2 <= 64'h0;
    end else if (io_clear) begin
      reg_file_2 <= 64'h0;
    end else if (write_en) begin
      if (2'h2 == write_addr[1:0]) begin
        if (io_instruction_valid) begin
          reg_file_2 <= _GEN_28[63:0];
        end else begin
          reg_file_2 <= 64'h0;
        end
      end
    end
    if (reset) begin
      reg_file_1 <= 64'h0;
    end else if (io_clear) begin
      reg_file_1 <= 64'h0;
    end else if (write_en) begin
      if (2'h1 == write_addr[1:0]) begin
        if (io_instruction_valid) begin
          reg_file_1 <= _GEN_28[63:0];
        end else begin
          reg_file_1 <= 64'h0;
        end
      end
    end
    if (reset) begin
      reg_file_0 <= 64'h0;
    end else if (io_clear) begin
      reg_file_0 <= 64'h0;
    end else if (write_en) begin
      if (2'h0 == write_addr[1:0]) begin
        if (io_instruction_valid) begin
          reg_file_0 <= _GEN_28[63:0];
        end else begin
          reg_file_0 <= 64'h0;
        end
      end
    end
  end
endmodule
module Mux3(
  input  [63:0] io_in_hardCoded,
  input  [63:0] io_in_data,
  input  [63:0] io_in_tbe,
  input  [1:0]  io_in_select,
  output        io_out_valid,
  output [63:0] io_out_bits
);
  wire  _T = io_in_select == 2'h3; // @[ComputationUtils.scala 27:24]
  wire  _T_1 = io_in_select == 2'h2; // @[ComputationUtils.scala 29:31]
  wire  _T_2 = io_in_select == 2'h1; // @[ComputationUtils.scala 31:31]
  wire [63:0] _GEN_0 = _T_2 ? io_in_tbe : 64'h0; // @[ComputationUtils.scala 31:40]
  wire [63:0] _GEN_1 = _T_1 ? io_in_data : _GEN_0; // @[ComputationUtils.scala 29:40]
  wire [63:0] result = _T ? io_in_hardCoded : _GEN_1; // @[ComputationUtils.scala 27:33]
  assign io_out_valid = result != 64'h0; // @[ComputationUtils.scala 38:18]
  assign io_out_bits = _T ? io_in_hardCoded : _GEN_1; // @[ComputationUtils.scala 37:17]
endmodule
module programmableCache(
  input         clock,
  input         reset,
  output        io_in_cpu_ready,
  input         io_in_cpu_valid,
  input  [1:0]  io_in_cpu_bits_event,
  input  [31:0] io_in_cpu_bits_addr,
  input  [63:0] io_in_cpu_bits_data,
  output        io_in_memCtrl_ready,
  input         io_in_memCtrl_valid,
  input  [1:0]  io_in_memCtrl_bits_event,
  input  [31:0] io_in_memCtrl_bits_addr,
  input  [63:0] io_in_memCtrl_bits_data,
  output        io_in_otherNodes_ready,
  input         io_in_otherNodes_valid,
  input  [1:0]  io_in_otherNodes_bits_event,
  input  [31:0] io_in_otherNodes_bits_addr,
  input  [63:0] io_in_otherNodes_bits_data,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_req_addr,
  output [7:0]  io_out_req_bits_req_inst,
  output [63:0] io_out_req_bits_req_data,
  output        io_out_resp_valid,
  output [31:0] io_out_resp_bits_addr,
  output        _T_814_0,
  output        _T_808_0,
  output        _T_819_0,
  output        hitLD_0,
  output        missLD_0,
  output        _T_811_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  cache_clock; // @[programmableCache.scala 52:26]
  wire  cache_reset; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_0_req_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_cpu_0_req_bits_addr; // @[programmableCache.scala 52:26]
  wire [27:0] cache_io_cpu_0_req_bits_command; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_0_req_bits_way; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_0_req_bits_replaceWay; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_0_resp_valid; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_0_resp_bits_iswrite; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_0_resp_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_1_req_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_cpu_1_req_bits_addr; // @[programmableCache.scala 52:26]
  wire [27:0] cache_io_cpu_1_req_bits_command; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_1_req_bits_way; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_1_req_bits_replaceWay; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_1_resp_valid; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_1_resp_bits_iswrite; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_1_resp_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_2_req_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_cpu_2_req_bits_addr; // @[programmableCache.scala 52:26]
  wire [27:0] cache_io_cpu_2_req_bits_command; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_2_req_bits_way; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_2_req_bits_replaceWay; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_2_resp_valid; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_2_resp_bits_iswrite; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_2_resp_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_3_req_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_cpu_3_req_bits_addr; // @[programmableCache.scala 52:26]
  wire [27:0] cache_io_cpu_3_req_bits_command; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_3_req_bits_way; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_3_req_bits_replaceWay; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_3_resp_valid; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_3_resp_bits_iswrite; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_3_resp_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_4_req_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_cpu_4_req_bits_addr; // @[programmableCache.scala 52:26]
  wire [27:0] cache_io_cpu_4_req_bits_command; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_4_req_bits_way; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_4_req_bits_replaceWay; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_4_resp_valid; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_4_resp_bits_iswrite; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_4_resp_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_5_req_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_cpu_5_req_bits_addr; // @[programmableCache.scala 52:26]
  wire [27:0] cache_io_cpu_5_req_bits_command; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_5_req_bits_way; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_5_req_bits_replaceWay; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_5_resp_valid; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_5_resp_bits_iswrite; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_5_resp_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_6_req_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_cpu_6_req_bits_addr; // @[programmableCache.scala 52:26]
  wire [27:0] cache_io_cpu_6_req_bits_command; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_6_req_bits_way; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_6_req_bits_replaceWay; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_6_resp_valid; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_6_resp_bits_iswrite; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_6_resp_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_7_req_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_cpu_7_req_bits_addr; // @[programmableCache.scala 52:26]
  wire [63:0] cache_io_cpu_7_req_bits_data; // @[programmableCache.scala 52:26]
  wire [27:0] cache_io_cpu_7_req_bits_command; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_7_req_bits_way; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_7_req_bits_replaceWay; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_7_resp_valid; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_7_resp_bits_iswrite; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_cpu_7_resp_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_probe_req_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_probe_req_bits_addr; // @[programmableCache.scala 52:26]
  wire [27:0] cache_io_probe_req_bits_command; // @[programmableCache.scala 52:26]
  wire  cache_io_probe_resp_valid; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_probe_resp_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_probe_multiWay_valid; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_probe_multiWay_bits_way_0; // @[programmableCache.scala 52:26]
  wire [1:0] cache_io_probe_multiWay_bits_way_1; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_probe_multiWay_bits_addr; // @[programmableCache.scala 52:26]
  wire  cache_io_bipassLD_in_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_bipassLD_in_bits_addr; // @[programmableCache.scala 52:26]
  wire [2:0] cache_io_bipassLD_in_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_bipassLD_out_valid; // @[programmableCache.scala 52:26]
  wire [63:0] cache_io_bipassLD_out_bits_data; // @[programmableCache.scala 52:26]
  wire  tbe_clock; // @[programmableCache.scala 53:26]
  wire  tbe_reset; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_0_valid; // @[programmableCache.scala 53:26]
  wire [63:0] tbe_io_write_0_bits_addr; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_0_bits_command; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_0_bits_mask; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_0_bits_inputTBE_state_state; // @[programmableCache.scala 53:26]
  wire [2:0] tbe_io_write_0_bits_inputTBE_way; // @[programmableCache.scala 53:26]
  wire [31:0] tbe_io_write_0_bits_inputTBE_fields_0; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_1_valid; // @[programmableCache.scala 53:26]
  wire [63:0] tbe_io_write_1_bits_addr; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_1_bits_command; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_1_bits_mask; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_1_bits_inputTBE_state_state; // @[programmableCache.scala 53:26]
  wire [2:0] tbe_io_write_1_bits_inputTBE_way; // @[programmableCache.scala 53:26]
  wire [31:0] tbe_io_write_1_bits_inputTBE_fields_0; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_2_valid; // @[programmableCache.scala 53:26]
  wire [63:0] tbe_io_write_2_bits_addr; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_2_bits_command; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_2_bits_mask; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_2_bits_inputTBE_state_state; // @[programmableCache.scala 53:26]
  wire [2:0] tbe_io_write_2_bits_inputTBE_way; // @[programmableCache.scala 53:26]
  wire [31:0] tbe_io_write_2_bits_inputTBE_fields_0; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_3_valid; // @[programmableCache.scala 53:26]
  wire [63:0] tbe_io_write_3_bits_addr; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_3_bits_command; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_3_bits_mask; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_3_bits_inputTBE_state_state; // @[programmableCache.scala 53:26]
  wire [2:0] tbe_io_write_3_bits_inputTBE_way; // @[programmableCache.scala 53:26]
  wire [31:0] tbe_io_write_3_bits_inputTBE_fields_0; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_4_valid; // @[programmableCache.scala 53:26]
  wire [63:0] tbe_io_write_4_bits_addr; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_4_bits_command; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_4_bits_mask; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_4_bits_inputTBE_state_state; // @[programmableCache.scala 53:26]
  wire [2:0] tbe_io_write_4_bits_inputTBE_way; // @[programmableCache.scala 53:26]
  wire [31:0] tbe_io_write_4_bits_inputTBE_fields_0; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_5_valid; // @[programmableCache.scala 53:26]
  wire [63:0] tbe_io_write_5_bits_addr; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_5_bits_command; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_5_bits_mask; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_5_bits_inputTBE_state_state; // @[programmableCache.scala 53:26]
  wire [2:0] tbe_io_write_5_bits_inputTBE_way; // @[programmableCache.scala 53:26]
  wire [31:0] tbe_io_write_5_bits_inputTBE_fields_0; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_6_valid; // @[programmableCache.scala 53:26]
  wire [63:0] tbe_io_write_6_bits_addr; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_6_bits_command; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_6_bits_mask; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_6_bits_inputTBE_state_state; // @[programmableCache.scala 53:26]
  wire [2:0] tbe_io_write_6_bits_inputTBE_way; // @[programmableCache.scala 53:26]
  wire [31:0] tbe_io_write_6_bits_inputTBE_fields_0; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_7_valid; // @[programmableCache.scala 53:26]
  wire [63:0] tbe_io_write_7_bits_addr; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_7_bits_command; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_7_bits_mask; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_7_bits_inputTBE_state_state; // @[programmableCache.scala 53:26]
  wire [2:0] tbe_io_write_7_bits_inputTBE_way; // @[programmableCache.scala 53:26]
  wire [31:0] tbe_io_write_7_bits_inputTBE_fields_0; // @[programmableCache.scala 53:26]
  wire  tbe_io_read_valid; // @[programmableCache.scala 53:26]
  wire [63:0] tbe_io_read_bits_addr; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_outputTBE_bits_state_state; // @[programmableCache.scala 53:26]
  wire [2:0] tbe_io_outputTBE_bits_way; // @[programmableCache.scala 53:26]
  wire [31:0] tbe_io_outputTBE_bits_fields_0; // @[programmableCache.scala 53:26]
  wire  tbe_io_isFull; // @[programmableCache.scala 53:26]
  wire  lockMem_clock; // @[programmableCache.scala 54:26]
  wire  lockMem_reset; // @[programmableCache.scala 54:26]
  wire  lockMem_io_lock_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_lock_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  lockMem_io_probe_out_valid; // @[programmableCache.scala 54:26]
  wire  lockMem_io_probe_out_bits; // @[programmableCache.scala 54:26]
  wire  lockMem_io_probe_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_probe_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  lockMem_io_unLock_0_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_unLock_0_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  lockMem_io_unLock_1_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_unLock_1_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  lockMem_io_unLock_2_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_unLock_2_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  lockMem_io_unLock_3_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_unLock_3_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  lockMem_io_unLock_4_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_unLock_4_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  lockMem_io_unLock_5_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_unLock_5_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  lockMem_io_unLock_6_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_unLock_6_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  lockMem_io_unLock_7_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_unLock_7_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  stateMem_clock; // @[programmableCache.scala 55:27]
  wire  stateMem_reset; // @[programmableCache.scala 55:27]
  wire  stateMem_io_in_0_valid; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_0_bits_state_state; // @[programmableCache.scala 55:27]
  wire [31:0] stateMem_io_in_0_bits_addr; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_0_bits_way; // @[programmableCache.scala 55:27]
  wire  stateMem_io_in_1_valid; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_1_bits_state_state; // @[programmableCache.scala 55:27]
  wire [31:0] stateMem_io_in_1_bits_addr; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_1_bits_way; // @[programmableCache.scala 55:27]
  wire  stateMem_io_in_2_valid; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_2_bits_state_state; // @[programmableCache.scala 55:27]
  wire [31:0] stateMem_io_in_2_bits_addr; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_2_bits_way; // @[programmableCache.scala 55:27]
  wire  stateMem_io_in_3_valid; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_3_bits_state_state; // @[programmableCache.scala 55:27]
  wire [31:0] stateMem_io_in_3_bits_addr; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_3_bits_way; // @[programmableCache.scala 55:27]
  wire  stateMem_io_in_4_valid; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_4_bits_state_state; // @[programmableCache.scala 55:27]
  wire [31:0] stateMem_io_in_4_bits_addr; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_4_bits_way; // @[programmableCache.scala 55:27]
  wire  stateMem_io_in_5_valid; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_5_bits_state_state; // @[programmableCache.scala 55:27]
  wire [31:0] stateMem_io_in_5_bits_addr; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_5_bits_way; // @[programmableCache.scala 55:27]
  wire  stateMem_io_in_6_valid; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_6_bits_state_state; // @[programmableCache.scala 55:27]
  wire [31:0] stateMem_io_in_6_bits_addr; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_6_bits_way; // @[programmableCache.scala 55:27]
  wire  stateMem_io_in_7_valid; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_7_bits_state_state; // @[programmableCache.scala 55:27]
  wire [31:0] stateMem_io_in_7_bits_addr; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_7_bits_way; // @[programmableCache.scala 55:27]
  wire  stateMem_io_in_8_valid; // @[programmableCache.scala 55:27]
  wire [31:0] stateMem_io_in_8_bits_addr; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_8_bits_way; // @[programmableCache.scala 55:27]
  wire  stateMem_io_out_valid; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_out_bits_state; // @[programmableCache.scala 55:27]
  wire  pc_clock; // @[programmableCache.scala 56:26]
  wire  pc_reset; // @[programmableCache.scala 56:26]
  wire  pc_io_write_ready; // @[programmableCache.scala 56:26]
  wire  pc_io_write_valid; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_write_bits_addr; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_write_bits_way; // @[programmableCache.scala 56:26]
  wire [63:0] pc_io_write_bits_data; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_write_bits_replaceWay; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_write_bits_tbeFields_0; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_write_bits_pc; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_0_in_bits_data_way; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_0_in_bits_data_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_0_in_bits_data_valid; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_0_out_bits_addr; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_0_out_bits_way; // @[programmableCache.scala 56:26]
  wire [63:0] pc_io_read_0_out_bits_data; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_0_out_bits_replaceWay; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_0_out_bits_tbeFields_0; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_0_out_bits_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_0_out_bits_valid; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_1_in_bits_data_way; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_1_in_bits_data_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_1_in_bits_data_valid; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_1_out_bits_addr; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_1_out_bits_way; // @[programmableCache.scala 56:26]
  wire [63:0] pc_io_read_1_out_bits_data; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_1_out_bits_replaceWay; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_1_out_bits_tbeFields_0; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_1_out_bits_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_1_out_bits_valid; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_2_in_bits_data_way; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_2_in_bits_data_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_2_in_bits_data_valid; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_2_out_bits_addr; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_2_out_bits_way; // @[programmableCache.scala 56:26]
  wire [63:0] pc_io_read_2_out_bits_data; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_2_out_bits_replaceWay; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_2_out_bits_tbeFields_0; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_2_out_bits_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_2_out_bits_valid; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_3_in_bits_data_way; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_3_in_bits_data_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_3_in_bits_data_valid; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_3_out_bits_addr; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_3_out_bits_way; // @[programmableCache.scala 56:26]
  wire [63:0] pc_io_read_3_out_bits_data; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_3_out_bits_replaceWay; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_3_out_bits_tbeFields_0; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_3_out_bits_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_3_out_bits_valid; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_4_in_bits_data_way; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_4_in_bits_data_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_4_in_bits_data_valid; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_4_out_bits_addr; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_4_out_bits_way; // @[programmableCache.scala 56:26]
  wire [63:0] pc_io_read_4_out_bits_data; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_4_out_bits_replaceWay; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_4_out_bits_tbeFields_0; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_4_out_bits_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_4_out_bits_valid; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_5_in_bits_data_way; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_5_in_bits_data_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_5_in_bits_data_valid; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_5_out_bits_addr; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_5_out_bits_way; // @[programmableCache.scala 56:26]
  wire [63:0] pc_io_read_5_out_bits_data; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_5_out_bits_replaceWay; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_5_out_bits_tbeFields_0; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_5_out_bits_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_5_out_bits_valid; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_6_in_bits_data_way; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_6_in_bits_data_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_6_in_bits_data_valid; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_6_out_bits_addr; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_6_out_bits_way; // @[programmableCache.scala 56:26]
  wire [63:0] pc_io_read_6_out_bits_data; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_6_out_bits_replaceWay; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_6_out_bits_tbeFields_0; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_6_out_bits_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_6_out_bits_valid; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_7_in_bits_data_way; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_7_in_bits_data_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_7_in_bits_data_valid; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_7_out_bits_addr; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_7_out_bits_way; // @[programmableCache.scala 56:26]
  wire [63:0] pc_io_read_7_out_bits_data; // @[programmableCache.scala 56:26]
  wire [1:0] pc_io_read_7_out_bits_replaceWay; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_7_out_bits_tbeFields_0; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_7_out_bits_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_7_out_bits_valid; // @[programmableCache.scala 56:26]
  wire  pc_io_isFull; // @[programmableCache.scala 56:26]
  wire  inputArbiter_io_in_0_valid; // @[programmableCache.scala 57:33]
  wire [1:0] inputArbiter_io_in_0_bits_event; // @[programmableCache.scala 57:33]
  wire [31:0] inputArbiter_io_in_0_bits_addr; // @[programmableCache.scala 57:33]
  wire [63:0] inputArbiter_io_in_0_bits_data; // @[programmableCache.scala 57:33]
  wire  inputArbiter_io_in_1_ready; // @[programmableCache.scala 57:33]
  wire  inputArbiter_io_in_1_valid; // @[programmableCache.scala 57:33]
  wire [1:0] inputArbiter_io_in_1_bits_event; // @[programmableCache.scala 57:33]
  wire [31:0] inputArbiter_io_in_1_bits_addr; // @[programmableCache.scala 57:33]
  wire [63:0] inputArbiter_io_in_1_bits_data; // @[programmableCache.scala 57:33]
  wire  inputArbiter_io_in_2_valid; // @[programmableCache.scala 57:33]
  wire [1:0] inputArbiter_io_in_2_bits_event; // @[programmableCache.scala 57:33]
  wire [31:0] inputArbiter_io_in_2_bits_addr; // @[programmableCache.scala 57:33]
  wire [63:0] inputArbiter_io_in_2_bits_data; // @[programmableCache.scala 57:33]
  wire  inputArbiter_io_in_3_valid; // @[programmableCache.scala 57:33]
  wire [1:0] inputArbiter_io_in_3_bits_event; // @[programmableCache.scala 57:33]
  wire [31:0] inputArbiter_io_in_3_bits_addr; // @[programmableCache.scala 57:33]
  wire [63:0] inputArbiter_io_in_3_bits_data; // @[programmableCache.scala 57:33]
  wire  inputArbiter_io_out_ready; // @[programmableCache.scala 57:33]
  wire  inputArbiter_io_out_valid; // @[programmableCache.scala 57:33]
  wire [1:0] inputArbiter_io_out_bits_event; // @[programmableCache.scala 57:33]
  wire [31:0] inputArbiter_io_out_bits_addr; // @[programmableCache.scala 57:33]
  wire [63:0] inputArbiter_io_out_bits_data; // @[programmableCache.scala 57:33]
  wire [1:0] inputArbiter_io_chosen; // @[programmableCache.scala 57:33]
  wire  outReqArbiter_clock; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_0_ready; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_0_valid; // @[programmableCache.scala 58:33]
  wire [31:0] outReqArbiter_io_in_0_bits_req_addr; // @[programmableCache.scala 58:33]
  wire [7:0] outReqArbiter_io_in_0_bits_req_inst; // @[programmableCache.scala 58:33]
  wire [63:0] outReqArbiter_io_in_0_bits_req_data; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_1_ready; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_1_valid; // @[programmableCache.scala 58:33]
  wire [31:0] outReqArbiter_io_in_1_bits_req_addr; // @[programmableCache.scala 58:33]
  wire [7:0] outReqArbiter_io_in_1_bits_req_inst; // @[programmableCache.scala 58:33]
  wire [63:0] outReqArbiter_io_in_1_bits_req_data; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_2_ready; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_2_valid; // @[programmableCache.scala 58:33]
  wire [31:0] outReqArbiter_io_in_2_bits_req_addr; // @[programmableCache.scala 58:33]
  wire [7:0] outReqArbiter_io_in_2_bits_req_inst; // @[programmableCache.scala 58:33]
  wire [63:0] outReqArbiter_io_in_2_bits_req_data; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_3_ready; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_3_valid; // @[programmableCache.scala 58:33]
  wire [31:0] outReqArbiter_io_in_3_bits_req_addr; // @[programmableCache.scala 58:33]
  wire [7:0] outReqArbiter_io_in_3_bits_req_inst; // @[programmableCache.scala 58:33]
  wire [63:0] outReqArbiter_io_in_3_bits_req_data; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_4_ready; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_4_valid; // @[programmableCache.scala 58:33]
  wire [31:0] outReqArbiter_io_in_4_bits_req_addr; // @[programmableCache.scala 58:33]
  wire [7:0] outReqArbiter_io_in_4_bits_req_inst; // @[programmableCache.scala 58:33]
  wire [63:0] outReqArbiter_io_in_4_bits_req_data; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_5_ready; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_5_valid; // @[programmableCache.scala 58:33]
  wire [31:0] outReqArbiter_io_in_5_bits_req_addr; // @[programmableCache.scala 58:33]
  wire [7:0] outReqArbiter_io_in_5_bits_req_inst; // @[programmableCache.scala 58:33]
  wire [63:0] outReqArbiter_io_in_5_bits_req_data; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_6_ready; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_6_valid; // @[programmableCache.scala 58:33]
  wire [31:0] outReqArbiter_io_in_6_bits_req_addr; // @[programmableCache.scala 58:33]
  wire [7:0] outReqArbiter_io_in_6_bits_req_inst; // @[programmableCache.scala 58:33]
  wire [63:0] outReqArbiter_io_in_6_bits_req_data; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_7_ready; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_in_7_valid; // @[programmableCache.scala 58:33]
  wire [31:0] outReqArbiter_io_in_7_bits_req_addr; // @[programmableCache.scala 58:33]
  wire [7:0] outReqArbiter_io_in_7_bits_req_inst; // @[programmableCache.scala 58:33]
  wire [63:0] outReqArbiter_io_in_7_bits_req_data; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_out_valid; // @[programmableCache.scala 58:33]
  wire [31:0] outReqArbiter_io_out_bits_req_addr; // @[programmableCache.scala 58:33]
  wire [7:0] outReqArbiter_io_out_bits_req_inst; // @[programmableCache.scala 58:33]
  wire [63:0] outReqArbiter_io_out_bits_req_data; // @[programmableCache.scala 58:33]
  wire [2:0] outReqArbiter_io_chosen; // @[programmableCache.scala 58:33]
  wire  outRespArbiter_io_in_0_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_in_0_bits_addr; // @[programmableCache.scala 59:33]
  wire  outRespArbiter_io_in_1_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_in_1_bits_addr; // @[programmableCache.scala 59:33]
  wire  outRespArbiter_io_in_2_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_in_2_bits_addr; // @[programmableCache.scala 59:33]
  wire  outRespArbiter_io_in_3_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_in_3_bits_addr; // @[programmableCache.scala 59:33]
  wire  outRespArbiter_io_in_4_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_in_4_bits_addr; // @[programmableCache.scala 59:33]
  wire  outRespArbiter_io_in_5_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_in_5_bits_addr; // @[programmableCache.scala 59:33]
  wire  outRespArbiter_io_in_6_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_in_6_bits_addr; // @[programmableCache.scala 59:33]
  wire  outRespArbiter_io_in_7_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_in_7_bits_addr; // @[programmableCache.scala 59:33]
  wire  outRespArbiter_io_in_8_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_in_8_bits_addr; // @[programmableCache.scala 59:33]
  wire  outRespArbiter_io_out_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_out_bits_addr; // @[programmableCache.scala 59:33]
  wire  feedbackArbiter_io_in_0_ready; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_0_valid; // @[programmableCache.scala 60:34]
  wire [1:0] feedbackArbiter_io_in_0_bits_event; // @[programmableCache.scala 60:34]
  wire [31:0] feedbackArbiter_io_in_0_bits_addr; // @[programmableCache.scala 60:34]
  wire [63:0] feedbackArbiter_io_in_0_bits_data; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_1_ready; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_1_valid; // @[programmableCache.scala 60:34]
  wire [1:0] feedbackArbiter_io_in_1_bits_event; // @[programmableCache.scala 60:34]
  wire [31:0] feedbackArbiter_io_in_1_bits_addr; // @[programmableCache.scala 60:34]
  wire [63:0] feedbackArbiter_io_in_1_bits_data; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_2_ready; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_2_valid; // @[programmableCache.scala 60:34]
  wire [1:0] feedbackArbiter_io_in_2_bits_event; // @[programmableCache.scala 60:34]
  wire [31:0] feedbackArbiter_io_in_2_bits_addr; // @[programmableCache.scala 60:34]
  wire [63:0] feedbackArbiter_io_in_2_bits_data; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_3_ready; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_3_valid; // @[programmableCache.scala 60:34]
  wire [1:0] feedbackArbiter_io_in_3_bits_event; // @[programmableCache.scala 60:34]
  wire [31:0] feedbackArbiter_io_in_3_bits_addr; // @[programmableCache.scala 60:34]
  wire [63:0] feedbackArbiter_io_in_3_bits_data; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_4_ready; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_4_valid; // @[programmableCache.scala 60:34]
  wire [1:0] feedbackArbiter_io_in_4_bits_event; // @[programmableCache.scala 60:34]
  wire [31:0] feedbackArbiter_io_in_4_bits_addr; // @[programmableCache.scala 60:34]
  wire [63:0] feedbackArbiter_io_in_4_bits_data; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_5_ready; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_5_valid; // @[programmableCache.scala 60:34]
  wire [1:0] feedbackArbiter_io_in_5_bits_event; // @[programmableCache.scala 60:34]
  wire [31:0] feedbackArbiter_io_in_5_bits_addr; // @[programmableCache.scala 60:34]
  wire [63:0] feedbackArbiter_io_in_5_bits_data; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_6_ready; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_6_valid; // @[programmableCache.scala 60:34]
  wire [1:0] feedbackArbiter_io_in_6_bits_event; // @[programmableCache.scala 60:34]
  wire [31:0] feedbackArbiter_io_in_6_bits_addr; // @[programmableCache.scala 60:34]
  wire [63:0] feedbackArbiter_io_in_6_bits_data; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_7_ready; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_7_valid; // @[programmableCache.scala 60:34]
  wire [1:0] feedbackArbiter_io_in_7_bits_event; // @[programmableCache.scala 60:34]
  wire [31:0] feedbackArbiter_io_in_7_bits_addr; // @[programmableCache.scala 60:34]
  wire [63:0] feedbackArbiter_io_in_7_bits_data; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_out_ready; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_out_valid; // @[programmableCache.scala 60:34]
  wire [1:0] feedbackArbiter_io_out_bits_event; // @[programmableCache.scala 60:34]
  wire [31:0] feedbackArbiter_io_out_bits_addr; // @[programmableCache.scala 60:34]
  wire [63:0] feedbackArbiter_io_out_bits_data; // @[programmableCache.scala 60:34]
  wire  input__clock; // @[programmableCache.scala 90:23]
  wire  input__reset; // @[programmableCache.scala 90:23]
  wire  input__io_enq_ready; // @[programmableCache.scala 90:23]
  wire  input__io_enq_valid; // @[programmableCache.scala 90:23]
  wire [1:0] input__io_enq_bits_inst_event; // @[programmableCache.scala 90:23]
  wire [31:0] input__io_enq_bits_inst_addr; // @[programmableCache.scala 90:23]
  wire [63:0] input__io_enq_bits_inst_data; // @[programmableCache.scala 90:23]
  wire [1:0] input__io_enq_bits_tbeOut_state_state; // @[programmableCache.scala 90:23]
  wire [2:0] input__io_enq_bits_tbeOut_way; // @[programmableCache.scala 90:23]
  wire [31:0] input__io_enq_bits_tbeOut_fields_0; // @[programmableCache.scala 90:23]
  wire  input__io_deq_ready; // @[programmableCache.scala 90:23]
  wire  input__io_deq_valid; // @[programmableCache.scala 90:23]
  wire [1:0] input__io_deq_bits_inst_event; // @[programmableCache.scala 90:23]
  wire [31:0] input__io_deq_bits_inst_addr; // @[programmableCache.scala 90:23]
  wire [63:0] input__io_deq_bits_inst_data; // @[programmableCache.scala 90:23]
  wire [1:0] input__io_deq_bits_tbeOut_state_state; // @[programmableCache.scala 90:23]
  wire [2:0] input__io_deq_bits_tbeOut_way; // @[programmableCache.scala 90:23]
  wire [31:0] input__io_deq_bits_tbeOut_fields_0; // @[programmableCache.scala 90:23]
  wire  respPortQueue_0_clock; // @[programmableCache.scala 93:27]
  wire  respPortQueue_0_reset; // @[programmableCache.scala 93:27]
  wire  respPortQueue_0_io_enq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_0_io_enq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_0_io_enq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_0_io_enq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_0_io_enq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_0_io_deq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_0_io_deq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_0_io_deq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_0_io_deq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_0_io_deq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_1_clock; // @[programmableCache.scala 93:27]
  wire  respPortQueue_1_reset; // @[programmableCache.scala 93:27]
  wire  respPortQueue_1_io_enq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_1_io_enq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_1_io_enq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_1_io_enq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_1_io_enq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_1_io_deq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_1_io_deq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_1_io_deq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_1_io_deq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_1_io_deq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_2_clock; // @[programmableCache.scala 93:27]
  wire  respPortQueue_2_reset; // @[programmableCache.scala 93:27]
  wire  respPortQueue_2_io_enq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_2_io_enq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_2_io_enq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_2_io_enq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_2_io_enq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_2_io_deq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_2_io_deq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_2_io_deq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_2_io_deq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_2_io_deq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_3_clock; // @[programmableCache.scala 93:27]
  wire  respPortQueue_3_reset; // @[programmableCache.scala 93:27]
  wire  respPortQueue_3_io_enq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_3_io_enq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_3_io_enq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_3_io_enq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_3_io_enq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_3_io_deq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_3_io_deq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_3_io_deq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_3_io_deq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_3_io_deq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_4_clock; // @[programmableCache.scala 93:27]
  wire  respPortQueue_4_reset; // @[programmableCache.scala 93:27]
  wire  respPortQueue_4_io_enq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_4_io_enq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_4_io_enq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_4_io_enq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_4_io_enq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_4_io_deq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_4_io_deq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_4_io_deq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_4_io_deq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_4_io_deq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_5_clock; // @[programmableCache.scala 93:27]
  wire  respPortQueue_5_reset; // @[programmableCache.scala 93:27]
  wire  respPortQueue_5_io_enq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_5_io_enq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_5_io_enq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_5_io_enq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_5_io_enq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_5_io_deq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_5_io_deq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_5_io_deq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_5_io_deq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_5_io_deq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_6_clock; // @[programmableCache.scala 93:27]
  wire  respPortQueue_6_reset; // @[programmableCache.scala 93:27]
  wire  respPortQueue_6_io_enq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_6_io_enq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_6_io_enq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_6_io_enq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_6_io_enq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_6_io_deq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_6_io_deq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_6_io_deq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_6_io_deq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_6_io_deq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_7_clock; // @[programmableCache.scala 93:27]
  wire  respPortQueue_7_reset; // @[programmableCache.scala 93:27]
  wire  respPortQueue_7_io_enq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_7_io_enq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_7_io_enq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_7_io_enq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_7_io_enq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_7_io_deq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_7_io_deq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_7_io_deq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_7_io_deq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_7_io_deq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_8_clock; // @[programmableCache.scala 93:27]
  wire  respPortQueue_8_reset; // @[programmableCache.scala 93:27]
  wire  respPortQueue_8_io_enq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_8_io_enq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_8_io_enq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_8_io_enq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_8_io_enq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_8_io_deq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_8_io_deq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_8_io_deq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_8_io_deq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_8_io_deq_bits_data; // @[programmableCache.scala 93:27]
  wire  reqPortQueue_0_clock; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_0_reset; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_0_io_enq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_0_io_enq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_0_io_enq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_0_io_enq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_0_io_enq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_0_io_deq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_0_io_deq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_0_io_deq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_0_io_deq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_0_io_deq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_1_clock; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_1_reset; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_1_io_enq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_1_io_enq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_1_io_enq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_1_io_enq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_1_io_enq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_1_io_deq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_1_io_deq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_1_io_deq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_1_io_deq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_1_io_deq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_2_clock; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_2_reset; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_2_io_enq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_2_io_enq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_2_io_enq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_2_io_enq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_2_io_enq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_2_io_deq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_2_io_deq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_2_io_deq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_2_io_deq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_2_io_deq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_3_clock; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_3_reset; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_3_io_enq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_3_io_enq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_3_io_enq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_3_io_enq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_3_io_enq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_3_io_deq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_3_io_deq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_3_io_deq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_3_io_deq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_3_io_deq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_4_clock; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_4_reset; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_4_io_enq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_4_io_enq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_4_io_enq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_4_io_enq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_4_io_enq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_4_io_deq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_4_io_deq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_4_io_deq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_4_io_deq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_4_io_deq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_5_clock; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_5_reset; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_5_io_enq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_5_io_enq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_5_io_enq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_5_io_enq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_5_io_enq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_5_io_deq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_5_io_deq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_5_io_deq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_5_io_deq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_5_io_deq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_6_clock; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_6_reset; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_6_io_enq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_6_io_enq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_6_io_enq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_6_io_enq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_6_io_enq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_6_io_deq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_6_io_deq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_6_io_deq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_6_io_deq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_6_io_deq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_7_clock; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_7_reset; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_7_io_enq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_7_io_enq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_7_io_enq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_7_io_enq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_7_io_enq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_7_io_deq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_7_io_deq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_7_io_deq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_7_io_deq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_7_io_deq_bits_data; // @[programmableCache.scala 98:27]
  wire  feedbackInQueue_0_clock; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_0_reset; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_0_io_enq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_0_io_enq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_0_io_enq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_0_io_enq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_0_io_enq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_0_io_deq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_0_io_deq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_0_io_deq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_0_io_deq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_0_io_deq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_1_clock; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_1_reset; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_1_io_enq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_1_io_enq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_1_io_enq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_1_io_enq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_1_io_enq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_1_io_deq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_1_io_deq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_1_io_deq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_1_io_deq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_1_io_deq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_2_clock; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_2_reset; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_2_io_enq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_2_io_enq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_2_io_enq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_2_io_enq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_2_io_enq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_2_io_deq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_2_io_deq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_2_io_deq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_2_io_deq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_2_io_deq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_3_clock; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_3_reset; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_3_io_enq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_3_io_enq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_3_io_enq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_3_io_enq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_3_io_enq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_3_io_deq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_3_io_deq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_3_io_deq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_3_io_deq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_3_io_deq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_4_clock; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_4_reset; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_4_io_enq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_4_io_enq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_4_io_enq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_4_io_enq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_4_io_enq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_4_io_deq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_4_io_deq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_4_io_deq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_4_io_deq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_4_io_deq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_5_clock; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_5_reset; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_5_io_enq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_5_io_enq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_5_io_enq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_5_io_enq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_5_io_enq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_5_io_deq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_5_io_deq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_5_io_deq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_5_io_deq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_5_io_deq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_6_clock; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_6_reset; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_6_io_enq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_6_io_enq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_6_io_enq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_6_io_enq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_6_io_enq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_6_io_deq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_6_io_deq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_6_io_deq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_6_io_deq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_6_io_deq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_7_clock; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_7_reset; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_7_io_enq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_7_io_enq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_7_io_enq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_7_io_enq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_7_io_enq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_7_io_deq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_7_io_deq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_7_io_deq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_7_io_deq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_7_io_deq_bits_data; // @[programmableCache.scala 104:27]
  wire  probeWay_clock; // @[programmableCache.scala 108:26]
  wire  probeWay_reset; // @[programmableCache.scala 108:26]
  wire  probeWay_io_enq_ready; // @[programmableCache.scala 108:26]
  wire  probeWay_io_enq_valid; // @[programmableCache.scala 108:26]
  wire [1:0] probeWay_io_enq_bits; // @[programmableCache.scala 108:26]
  wire  probeWay_io_deq_ready; // @[programmableCache.scala 108:26]
  wire  probeWay_io_deq_valid; // @[programmableCache.scala 108:26]
  wire [1:0] probeWay_io_deq_bits; // @[programmableCache.scala 108:26]
  wire  feedbackOutQueue_clock; // @[programmableCache.scala 165:34]
  wire  feedbackOutQueue_reset; // @[programmableCache.scala 165:34]
  wire  feedbackOutQueue_io_enq_ready; // @[programmableCache.scala 165:34]
  wire  feedbackOutQueue_io_enq_valid; // @[programmableCache.scala 165:34]
  wire [1:0] feedbackOutQueue_io_enq_bits_event; // @[programmableCache.scala 165:34]
  wire [31:0] feedbackOutQueue_io_enq_bits_addr; // @[programmableCache.scala 165:34]
  wire [63:0] feedbackOutQueue_io_enq_bits_data; // @[programmableCache.scala 165:34]
  wire  feedbackOutQueue_io_deq_ready; // @[programmableCache.scala 165:34]
  wire  feedbackOutQueue_io_deq_valid; // @[programmableCache.scala 165:34]
  wire [1:0] feedbackOutQueue_io_deq_bits_event; // @[programmableCache.scala 165:34]
  wire [31:0] feedbackOutQueue_io_deq_bits_addr; // @[programmableCache.scala 165:34]
  wire [63:0] feedbackOutQueue_io_deq_bits_data; // @[programmableCache.scala 165:34]
  wire  routineQueue_clock; // @[programmableCache.scala 166:30]
  wire  routineQueue_reset; // @[programmableCache.scala 166:30]
  wire  routineQueue_io_enq_ready; // @[programmableCache.scala 166:30]
  wire  routineQueue_io_enq_valid; // @[programmableCache.scala 166:30]
  wire [15:0] routineQueue_io_enq_bits; // @[programmableCache.scala 166:30]
  wire  routineQueue_io_deq_ready; // @[programmableCache.scala 166:30]
  wire  routineQueue_io_deq_valid; // @[programmableCache.scala 166:30]
  wire [15:0] routineQueue_io_deq_bits; // @[programmableCache.scala 166:30]
  wire  actionReg_0_clock; // @[programmableCache.scala 169:32]
  wire  actionReg_0_reset; // @[programmableCache.scala 169:32]
  wire  actionReg_0_io_enq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_0_io_enq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_0_io_enq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_0_io_enq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_0_io_enq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_0_io_enq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_0_io_enq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_0_io_enq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_0_io_enq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_0_io_deq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_0_io_deq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_0_io_deq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_0_io_deq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_0_io_deq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_0_io_deq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_0_io_deq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_0_io_deq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_0_io_deq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_1_clock; // @[programmableCache.scala 169:32]
  wire  actionReg_1_reset; // @[programmableCache.scala 169:32]
  wire  actionReg_1_io_enq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_1_io_enq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_1_io_enq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_1_io_enq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_1_io_enq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_1_io_enq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_1_io_enq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_1_io_enq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_1_io_enq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_1_io_deq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_1_io_deq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_1_io_deq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_1_io_deq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_1_io_deq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_1_io_deq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_1_io_deq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_1_io_deq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_1_io_deq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_2_clock; // @[programmableCache.scala 169:32]
  wire  actionReg_2_reset; // @[programmableCache.scala 169:32]
  wire  actionReg_2_io_enq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_2_io_enq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_2_io_enq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_2_io_enq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_2_io_enq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_2_io_enq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_2_io_enq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_2_io_enq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_2_io_enq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_2_io_deq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_2_io_deq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_2_io_deq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_2_io_deq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_2_io_deq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_2_io_deq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_2_io_deq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_2_io_deq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_2_io_deq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_3_clock; // @[programmableCache.scala 169:32]
  wire  actionReg_3_reset; // @[programmableCache.scala 169:32]
  wire  actionReg_3_io_enq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_3_io_enq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_3_io_enq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_3_io_enq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_3_io_enq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_3_io_enq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_3_io_enq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_3_io_enq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_3_io_enq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_3_io_deq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_3_io_deq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_3_io_deq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_3_io_deq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_3_io_deq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_3_io_deq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_3_io_deq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_3_io_deq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_3_io_deq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_4_clock; // @[programmableCache.scala 169:32]
  wire  actionReg_4_reset; // @[programmableCache.scala 169:32]
  wire  actionReg_4_io_enq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_4_io_enq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_4_io_enq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_4_io_enq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_4_io_enq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_4_io_enq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_4_io_enq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_4_io_enq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_4_io_enq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_4_io_deq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_4_io_deq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_4_io_deq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_4_io_deq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_4_io_deq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_4_io_deq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_4_io_deq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_4_io_deq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_4_io_deq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_5_clock; // @[programmableCache.scala 169:32]
  wire  actionReg_5_reset; // @[programmableCache.scala 169:32]
  wire  actionReg_5_io_enq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_5_io_enq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_5_io_enq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_5_io_enq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_5_io_enq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_5_io_enq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_5_io_enq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_5_io_enq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_5_io_enq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_5_io_deq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_5_io_deq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_5_io_deq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_5_io_deq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_5_io_deq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_5_io_deq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_5_io_deq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_5_io_deq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_5_io_deq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_6_clock; // @[programmableCache.scala 169:32]
  wire  actionReg_6_reset; // @[programmableCache.scala 169:32]
  wire  actionReg_6_io_enq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_6_io_enq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_6_io_enq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_6_io_enq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_6_io_enq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_6_io_enq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_6_io_enq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_6_io_enq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_6_io_enq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_6_io_deq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_6_io_deq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_6_io_deq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_6_io_deq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_6_io_deq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_6_io_deq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_6_io_deq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_6_io_deq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_6_io_deq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_7_clock; // @[programmableCache.scala 169:32]
  wire  actionReg_7_reset; // @[programmableCache.scala 169:32]
  wire  actionReg_7_io_enq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_7_io_enq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_7_io_enq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_7_io_enq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_7_io_enq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_7_io_enq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_7_io_enq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_7_io_enq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_7_io_enq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_7_io_deq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_7_io_deq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_7_io_deq_bits_addr; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_7_io_deq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_7_io_deq_bits_data; // @[programmableCache.scala 169:32]
  wire [1:0] actionReg_7_io_deq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_7_io_deq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_7_io_deq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_7_io_deq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  mimoQ_clock; // @[programmableCache.scala 173:24]
  wire  mimoQ_reset; // @[programmableCache.scala 173:24]
  wire  mimoQ_io_enq_ready; // @[programmableCache.scala 173:24]
  wire  mimoQ_io_enq_valid; // @[programmableCache.scala 173:24]
  wire [1:0] mimoQ_io_enq_bits_0_way; // @[programmableCache.scala 173:24]
  wire [31:0] mimoQ_io_enq_bits_0_addr; // @[programmableCache.scala 173:24]
  wire [1:0] mimoQ_io_enq_bits_1_way; // @[programmableCache.scala 173:24]
  wire [31:0] mimoQ_io_enq_bits_1_addr; // @[programmableCache.scala 173:24]
  wire  mimoQ_io_deq_valid; // @[programmableCache.scala 173:24]
  wire [1:0] mimoQ_io_deq_bits_0_way; // @[programmableCache.scala 173:24]
  wire [31:0] mimoQ_io_deq_bits_0_addr; // @[programmableCache.scala 173:24]
  wire [3:0] mimoQ_io_count; // @[programmableCache.scala 173:24]
  wire  compUnit_0_clock; // @[programmableCache.scala 177:27]
  wire  compUnit_0_reset; // @[programmableCache.scala 177:27]
  wire  compUnit_0_io_instruction_valid; // @[programmableCache.scala 177:27]
  wire [27:0] compUnit_0_io_instruction_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_0_io_clear; // @[programmableCache.scala 177:27]
  wire  compUnit_0_io_op1_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_0_io_op1_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_0_io_op2_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_0_io_op2_bits; // @[programmableCache.scala 177:27]
  wire [15:0] compUnit_0_io_pc; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_0_io_reg_file_0; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_0_io_reg_file_1; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_0_io_reg_file_2; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_0_io_reg_file_3; // @[programmableCache.scala 177:27]
  wire  compUnit_1_clock; // @[programmableCache.scala 177:27]
  wire  compUnit_1_reset; // @[programmableCache.scala 177:27]
  wire  compUnit_1_io_instruction_valid; // @[programmableCache.scala 177:27]
  wire [27:0] compUnit_1_io_instruction_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_1_io_clear; // @[programmableCache.scala 177:27]
  wire  compUnit_1_io_op1_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_1_io_op1_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_1_io_op2_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_1_io_op2_bits; // @[programmableCache.scala 177:27]
  wire [15:0] compUnit_1_io_pc; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_1_io_reg_file_0; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_1_io_reg_file_1; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_1_io_reg_file_2; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_1_io_reg_file_3; // @[programmableCache.scala 177:27]
  wire  compUnit_2_clock; // @[programmableCache.scala 177:27]
  wire  compUnit_2_reset; // @[programmableCache.scala 177:27]
  wire  compUnit_2_io_instruction_valid; // @[programmableCache.scala 177:27]
  wire [27:0] compUnit_2_io_instruction_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_2_io_clear; // @[programmableCache.scala 177:27]
  wire  compUnit_2_io_op1_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_2_io_op1_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_2_io_op2_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_2_io_op2_bits; // @[programmableCache.scala 177:27]
  wire [15:0] compUnit_2_io_pc; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_2_io_reg_file_0; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_2_io_reg_file_1; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_2_io_reg_file_2; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_2_io_reg_file_3; // @[programmableCache.scala 177:27]
  wire  compUnit_3_clock; // @[programmableCache.scala 177:27]
  wire  compUnit_3_reset; // @[programmableCache.scala 177:27]
  wire  compUnit_3_io_instruction_valid; // @[programmableCache.scala 177:27]
  wire [27:0] compUnit_3_io_instruction_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_3_io_clear; // @[programmableCache.scala 177:27]
  wire  compUnit_3_io_op1_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_3_io_op1_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_3_io_op2_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_3_io_op2_bits; // @[programmableCache.scala 177:27]
  wire [15:0] compUnit_3_io_pc; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_3_io_reg_file_0; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_3_io_reg_file_1; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_3_io_reg_file_2; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_3_io_reg_file_3; // @[programmableCache.scala 177:27]
  wire  compUnit_4_clock; // @[programmableCache.scala 177:27]
  wire  compUnit_4_reset; // @[programmableCache.scala 177:27]
  wire  compUnit_4_io_instruction_valid; // @[programmableCache.scala 177:27]
  wire [27:0] compUnit_4_io_instruction_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_4_io_clear; // @[programmableCache.scala 177:27]
  wire  compUnit_4_io_op1_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_4_io_op1_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_4_io_op2_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_4_io_op2_bits; // @[programmableCache.scala 177:27]
  wire [15:0] compUnit_4_io_pc; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_4_io_reg_file_0; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_4_io_reg_file_1; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_4_io_reg_file_2; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_4_io_reg_file_3; // @[programmableCache.scala 177:27]
  wire  compUnit_5_clock; // @[programmableCache.scala 177:27]
  wire  compUnit_5_reset; // @[programmableCache.scala 177:27]
  wire  compUnit_5_io_instruction_valid; // @[programmableCache.scala 177:27]
  wire [27:0] compUnit_5_io_instruction_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_5_io_clear; // @[programmableCache.scala 177:27]
  wire  compUnit_5_io_op1_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_5_io_op1_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_5_io_op2_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_5_io_op2_bits; // @[programmableCache.scala 177:27]
  wire [15:0] compUnit_5_io_pc; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_5_io_reg_file_0; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_5_io_reg_file_1; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_5_io_reg_file_2; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_5_io_reg_file_3; // @[programmableCache.scala 177:27]
  wire  compUnit_6_clock; // @[programmableCache.scala 177:27]
  wire  compUnit_6_reset; // @[programmableCache.scala 177:27]
  wire  compUnit_6_io_instruction_valid; // @[programmableCache.scala 177:27]
  wire [27:0] compUnit_6_io_instruction_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_6_io_clear; // @[programmableCache.scala 177:27]
  wire  compUnit_6_io_op1_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_6_io_op1_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_6_io_op2_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_6_io_op2_bits; // @[programmableCache.scala 177:27]
  wire [15:0] compUnit_6_io_pc; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_6_io_reg_file_0; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_6_io_reg_file_1; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_6_io_reg_file_2; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_6_io_reg_file_3; // @[programmableCache.scala 177:27]
  wire  compUnit_7_clock; // @[programmableCache.scala 177:27]
  wire  compUnit_7_reset; // @[programmableCache.scala 177:27]
  wire  compUnit_7_io_instruction_valid; // @[programmableCache.scala 177:27]
  wire [27:0] compUnit_7_io_instruction_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_7_io_clear; // @[programmableCache.scala 177:27]
  wire  compUnit_7_io_op1_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_7_io_op1_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_7_io_op2_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_7_io_op2_bits; // @[programmableCache.scala 177:27]
  wire [15:0] compUnit_7_io_pc; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_7_io_reg_file_0; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_7_io_reg_file_1; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_7_io_reg_file_2; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_7_io_reg_file_3; // @[programmableCache.scala 177:27]
  wire [63:0] compUnitInput1_0_io_in_hardCoded; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_0_io_in_data; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_0_io_in_tbe; // @[programmableCache.scala 182:30]
  wire [1:0] compUnitInput1_0_io_in_select; // @[programmableCache.scala 182:30]
  wire  compUnitInput1_0_io_out_valid; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_0_io_out_bits; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_1_io_in_hardCoded; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_1_io_in_data; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_1_io_in_tbe; // @[programmableCache.scala 182:30]
  wire [1:0] compUnitInput1_1_io_in_select; // @[programmableCache.scala 182:30]
  wire  compUnitInput1_1_io_out_valid; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_1_io_out_bits; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_2_io_in_hardCoded; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_2_io_in_data; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_2_io_in_tbe; // @[programmableCache.scala 182:30]
  wire [1:0] compUnitInput1_2_io_in_select; // @[programmableCache.scala 182:30]
  wire  compUnitInput1_2_io_out_valid; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_2_io_out_bits; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_3_io_in_hardCoded; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_3_io_in_data; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_3_io_in_tbe; // @[programmableCache.scala 182:30]
  wire [1:0] compUnitInput1_3_io_in_select; // @[programmableCache.scala 182:30]
  wire  compUnitInput1_3_io_out_valid; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_3_io_out_bits; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_4_io_in_hardCoded; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_4_io_in_data; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_4_io_in_tbe; // @[programmableCache.scala 182:30]
  wire [1:0] compUnitInput1_4_io_in_select; // @[programmableCache.scala 182:30]
  wire  compUnitInput1_4_io_out_valid; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_4_io_out_bits; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_5_io_in_hardCoded; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_5_io_in_data; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_5_io_in_tbe; // @[programmableCache.scala 182:30]
  wire [1:0] compUnitInput1_5_io_in_select; // @[programmableCache.scala 182:30]
  wire  compUnitInput1_5_io_out_valid; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_5_io_out_bits; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_6_io_in_hardCoded; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_6_io_in_data; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_6_io_in_tbe; // @[programmableCache.scala 182:30]
  wire [1:0] compUnitInput1_6_io_in_select; // @[programmableCache.scala 182:30]
  wire  compUnitInput1_6_io_out_valid; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_6_io_out_bits; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_7_io_in_hardCoded; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_7_io_in_data; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_7_io_in_tbe; // @[programmableCache.scala 182:30]
  wire [1:0] compUnitInput1_7_io_in_select; // @[programmableCache.scala 182:30]
  wire  compUnitInput1_7_io_out_valid; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_7_io_out_bits; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput2_0_io_in_hardCoded; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_0_io_in_data; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_0_io_in_tbe; // @[programmableCache.scala 188:30]
  wire [1:0] compUnitInput2_0_io_in_select; // @[programmableCache.scala 188:30]
  wire  compUnitInput2_0_io_out_valid; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_0_io_out_bits; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_1_io_in_hardCoded; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_1_io_in_data; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_1_io_in_tbe; // @[programmableCache.scala 188:30]
  wire [1:0] compUnitInput2_1_io_in_select; // @[programmableCache.scala 188:30]
  wire  compUnitInput2_1_io_out_valid; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_1_io_out_bits; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_2_io_in_hardCoded; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_2_io_in_data; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_2_io_in_tbe; // @[programmableCache.scala 188:30]
  wire [1:0] compUnitInput2_2_io_in_select; // @[programmableCache.scala 188:30]
  wire  compUnitInput2_2_io_out_valid; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_2_io_out_bits; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_3_io_in_hardCoded; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_3_io_in_data; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_3_io_in_tbe; // @[programmableCache.scala 188:30]
  wire [1:0] compUnitInput2_3_io_in_select; // @[programmableCache.scala 188:30]
  wire  compUnitInput2_3_io_out_valid; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_3_io_out_bits; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_4_io_in_hardCoded; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_4_io_in_data; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_4_io_in_tbe; // @[programmableCache.scala 188:30]
  wire [1:0] compUnitInput2_4_io_in_select; // @[programmableCache.scala 188:30]
  wire  compUnitInput2_4_io_out_valid; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_4_io_out_bits; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_5_io_in_hardCoded; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_5_io_in_data; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_5_io_in_tbe; // @[programmableCache.scala 188:30]
  wire [1:0] compUnitInput2_5_io_in_select; // @[programmableCache.scala 188:30]
  wire  compUnitInput2_5_io_out_valid; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_5_io_out_bits; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_6_io_in_hardCoded; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_6_io_in_data; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_6_io_in_tbe; // @[programmableCache.scala 188:30]
  wire [1:0] compUnitInput2_6_io_in_select; // @[programmableCache.scala 188:30]
  wire  compUnitInput2_6_io_out_valid; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_6_io_out_bits; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_7_io_in_hardCoded; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_7_io_in_data; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_7_io_in_tbe; // @[programmableCache.scala 188:30]
  wire [1:0] compUnitInput2_7_io_in_select; // @[programmableCache.scala 188:30]
  wire  compUnitInput2_7_io_out_valid; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_7_io_out_bits; // @[programmableCache.scala 188:30]
  wire  _T_182 = input__io_deq_bits_tbeOut_state_state != 2'h0; // @[programmableCache.scala 293:55]
  wire [1:0] _T_183 = stateMem_io_out_valid ? stateMem_io_out_bits_state : 2'h0; // @[programmableCache.scala 293:120]
  wire [1:0] state = _T_182 ? input__io_deq_bits_tbeOut_state_state : _T_183; // @[programmableCache.scala 293:17]
  wire [3:0] routine = {input__io_deq_bits_inst_event,state}; // @[Cat.scala 29:58]
  reg  instUsed; // @[programmableCache.scala 197:27]
  reg  replStateReg_0; // @[programmableCache.scala 204:31]
  reg  replStateReg_1; // @[programmableCache.scala 204:31]
  wire [31:0] _GEN_1510 = {{24'd0}, actionReg_0_io_deq_bits_action_signals[7:0]}; // @[programmableCache.scala 247:78]
  wire [63:0] _GEN_1511 = {{60'd0}, actionReg_0_io_deq_bits_action_signals[11:8]}; // @[programmableCache.scala 249:78]
  wire [31:0] _GEN_1512 = {{24'd0}, actionReg_1_io_deq_bits_action_signals[7:0]}; // @[programmableCache.scala 247:78]
  wire [63:0] _GEN_1513 = {{60'd0}, actionReg_1_io_deq_bits_action_signals[11:8]}; // @[programmableCache.scala 249:78]
  wire [31:0] _GEN_1514 = {{24'd0}, actionReg_2_io_deq_bits_action_signals[7:0]}; // @[programmableCache.scala 247:78]
  wire [63:0] _GEN_1515 = {{60'd0}, actionReg_2_io_deq_bits_action_signals[11:8]}; // @[programmableCache.scala 249:78]
  wire [31:0] _GEN_1516 = {{24'd0}, actionReg_3_io_deq_bits_action_signals[7:0]}; // @[programmableCache.scala 247:78]
  wire [63:0] _GEN_1517 = {{60'd0}, actionReg_3_io_deq_bits_action_signals[11:8]}; // @[programmableCache.scala 249:78]
  wire [31:0] _GEN_1518 = {{24'd0}, actionReg_4_io_deq_bits_action_signals[7:0]}; // @[programmableCache.scala 247:78]
  wire [63:0] _GEN_1519 = {{60'd0}, actionReg_4_io_deq_bits_action_signals[11:8]}; // @[programmableCache.scala 249:78]
  wire [31:0] _GEN_1520 = {{24'd0}, actionReg_5_io_deq_bits_action_signals[7:0]}; // @[programmableCache.scala 247:78]
  wire [63:0] _GEN_1521 = {{60'd0}, actionReg_5_io_deq_bits_action_signals[11:8]}; // @[programmableCache.scala 249:78]
  wire [31:0] _GEN_1522 = {{24'd0}, actionReg_6_io_deq_bits_action_signals[7:0]}; // @[programmableCache.scala 247:78]
  wire [63:0] _GEN_1523 = {{60'd0}, actionReg_6_io_deq_bits_action_signals[11:8]}; // @[programmableCache.scala 249:78]
  wire [31:0] _GEN_1524 = {{24'd0}, actionReg_7_io_deq_bits_action_signals[7:0]}; // @[programmableCache.scala 247:78]
  wire [63:0] _GEN_1525 = {{60'd0}, actionReg_7_io_deq_bits_action_signals[11:8]}; // @[programmableCache.scala 249:78]
  wire  isLocked = lockMem_io_probe_out_valid & lockMem_io_probe_out_bits; // @[programmableCache.scala 323:21]
  wire  stallInput = isLocked | tbe_io_isFull; // @[programmableCache.scala 260:28]
  wire  hitEvent = 2'h0 == input__io_deq_bits_inst_event; // @[programmableCache.scala 264:35]
  wire  _T_171 = ~tbe_io_isFull; // @[programmableCache.scala 284:48]
  wire  _T_172 = input__io_enq_ready & _T_171; // @[programmableCache.scala 284:45]
  wire  _T_173 = ~stallInput; // @[programmableCache.scala 284:66]
  wire  instruction_ready = _T_172 & _T_173; // @[programmableCache.scala 284:63]
  wire  instruction_valid = inputArbiter_io_out_valid; // @[programmableCache.scala 110:27 programmableCache.scala 252:17]
  wire  _T_141 = instruction_ready & instruction_valid; // @[Decoupled.scala 40:37]
  wire [1:0] instruction_bits_event = inputArbiter_io_out_bits_event; // @[programmableCache.scala 110:27 programmableCache.scala 252:17]
  wire  _T_142 = 2'h0 == instruction_bits_event; // @[programmableCache.scala 267:59]
  wire  probeStart = _T_141 & _T_142; // @[programmableCache.scala 267:38]
  wire  getState = input__io_deq_ready & input__io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_149 = probeWay_io_deq_bits != 2'h2; // @[programmableCache.scala 275:46]
  wire  _T_150 = getState & _T_149; // @[programmableCache.scala 275:21]
  wire  _T_151 = stateMem_io_out_bits_state == 2'h3; // @[programmableCache.scala 275:90]
  wire  hit = _T_150 & _T_151; // @[programmableCache.scala 275:59]
  wire  _T_153 = hit & hitEvent; // @[programmableCache.scala 276:20]
  wire  _T_154 = getState & hitEvent; // @[programmableCache.scala 277:24]
  wire  _T_155 = stateMem_io_out_bits_state == 2'h0; // @[programmableCache.scala 277:71]
  wire  _T_156 = _T_154 & _T_155; // @[programmableCache.scala 277:39]
  wire  _T_158 = inputArbiter_io_chosen == 2'h0; // @[programmableCache.scala 279:77]
  wire  _T_159 = _T_141 & _T_158; // @[programmableCache.scala 279:51]
  wire  _T_161 = inputArbiter_io_chosen == 2'h3; // @[programmableCache.scala 280:76]
  wire  _T_162 = _T_141 & _T_161; // @[programmableCache.scala 280:50]
  wire  _T_164 = inputArbiter_io_chosen == 2'h2; // @[programmableCache.scala 281:77]
  wire  _T_167 = ~_T_141; // @[programmableCache.scala 283:20]
  wire  _T_168 = input__io_enq_ready & input__io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_169 = _T_168 | instUsed; // @[programmableCache.scala 283:63]
  wire  _T_170 = _T_167 & _T_169; // @[programmableCache.scala 283:40]
  wire  _T_175 = ~instUsed; // @[programmableCache.scala 286:48]
  wire  _T_176 = instruction_valid & _T_175; // @[programmableCache.scala 286:45]
  wire  _T_178 = _T_176 & _T_171; // @[programmableCache.scala 286:58]
  wire  maskField_0 = actionReg_0_io_deq_bits_action_signals[2]; // @[Gem5CacheLogic.scala 114:54]
  wire  _T_185 = ~maskField_0; // @[programmableCache.scala 303:84]
  wire [63:0] _GEN_207 = compUnit_0_io_reg_file_0; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_208 = 2'h1 == actionReg_0_io_deq_bits_action_signals[4:3] ? compUnit_0_io_reg_file_1 : _GEN_207; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_209 = 2'h2 == actionReg_0_io_deq_bits_action_signals[4:3] ? compUnit_0_io_reg_file_2 : _GEN_208; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_210 = 2'h3 == actionReg_0_io_deq_bits_action_signals[4:3] ? compUnit_0_io_reg_file_3 : _GEN_209; // @[programmableCache.scala 417:31]
  wire [31:0] tbeFieldUpdateSrc_0 = _GEN_210[31:0]; // @[programmableCache.scala 138:33 programmableCache.scala 417:31]
  wire  _T_280 = actionReg_0_io_deq_bits_action_actionType == 4'h3; // @[programmableCache.scala 373:73]
  wire  isStateAction_0 = _T_280 & actionReg_0_io_deq_valid; // @[programmableCache.scala 373:82]
  wire [1:0] tbeAction_0 = actionReg_0_io_deq_bits_action_signals[1:0]; // @[Gem5CacheLogic.scala 115:54]
  wire  _T_274 = actionReg_0_io_deq_bits_action_actionType == 4'h1; // @[programmableCache.scala 370:73]
  wire  isTBEAction_0 = _T_274 & actionReg_0_io_deq_valid; // @[programmableCache.scala 370:82]
  wire  maskField_1 = actionReg_1_io_deq_bits_action_signals[2]; // @[Gem5CacheLogic.scala 114:54]
  wire  _T_191 = ~maskField_1; // @[programmableCache.scala 303:84]
  wire [63:0] _GEN_388 = compUnit_1_io_reg_file_0; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_389 = 2'h1 == actionReg_1_io_deq_bits_action_signals[4:3] ? compUnit_1_io_reg_file_1 : _GEN_388; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_390 = 2'h2 == actionReg_1_io_deq_bits_action_signals[4:3] ? compUnit_1_io_reg_file_2 : _GEN_389; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_391 = 2'h3 == actionReg_1_io_deq_bits_action_signals[4:3] ? compUnit_1_io_reg_file_3 : _GEN_390; // @[programmableCache.scala 417:31]
  wire [31:0] tbeFieldUpdateSrc_1 = _GEN_391[31:0]; // @[programmableCache.scala 138:33 programmableCache.scala 417:31]
  wire  _T_337 = actionReg_1_io_deq_bits_action_actionType == 4'h3; // @[programmableCache.scala 373:73]
  wire  isStateAction_1 = _T_337 & actionReg_1_io_deq_valid; // @[programmableCache.scala 373:82]
  wire [1:0] tbeAction_1 = actionReg_1_io_deq_bits_action_signals[1:0]; // @[Gem5CacheLogic.scala 115:54]
  wire  _T_331 = actionReg_1_io_deq_bits_action_actionType == 4'h1; // @[programmableCache.scala 370:73]
  wire  isTBEAction_1 = _T_331 & actionReg_1_io_deq_valid; // @[programmableCache.scala 370:82]
  wire  maskField_2 = actionReg_2_io_deq_bits_action_signals[2]; // @[Gem5CacheLogic.scala 114:54]
  wire  _T_197 = ~maskField_2; // @[programmableCache.scala 303:84]
  wire [63:0] _GEN_569 = compUnit_2_io_reg_file_0; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_570 = 2'h1 == actionReg_2_io_deq_bits_action_signals[4:3] ? compUnit_2_io_reg_file_1 : _GEN_569; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_571 = 2'h2 == actionReg_2_io_deq_bits_action_signals[4:3] ? compUnit_2_io_reg_file_2 : _GEN_570; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_572 = 2'h3 == actionReg_2_io_deq_bits_action_signals[4:3] ? compUnit_2_io_reg_file_3 : _GEN_571; // @[programmableCache.scala 417:31]
  wire [31:0] tbeFieldUpdateSrc_2 = _GEN_572[31:0]; // @[programmableCache.scala 138:33 programmableCache.scala 417:31]
  wire  _T_394 = actionReg_2_io_deq_bits_action_actionType == 4'h3; // @[programmableCache.scala 373:73]
  wire  isStateAction_2 = _T_394 & actionReg_2_io_deq_valid; // @[programmableCache.scala 373:82]
  wire [1:0] tbeAction_2 = actionReg_2_io_deq_bits_action_signals[1:0]; // @[Gem5CacheLogic.scala 115:54]
  wire  _T_388 = actionReg_2_io_deq_bits_action_actionType == 4'h1; // @[programmableCache.scala 370:73]
  wire  isTBEAction_2 = _T_388 & actionReg_2_io_deq_valid; // @[programmableCache.scala 370:82]
  wire  maskField_3 = actionReg_3_io_deq_bits_action_signals[2]; // @[Gem5CacheLogic.scala 114:54]
  wire  _T_203 = ~maskField_3; // @[programmableCache.scala 303:84]
  wire [63:0] _GEN_750 = compUnit_3_io_reg_file_0; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_751 = 2'h1 == actionReg_3_io_deq_bits_action_signals[4:3] ? compUnit_3_io_reg_file_1 : _GEN_750; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_752 = 2'h2 == actionReg_3_io_deq_bits_action_signals[4:3] ? compUnit_3_io_reg_file_2 : _GEN_751; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_753 = 2'h3 == actionReg_3_io_deq_bits_action_signals[4:3] ? compUnit_3_io_reg_file_3 : _GEN_752; // @[programmableCache.scala 417:31]
  wire [31:0] tbeFieldUpdateSrc_3 = _GEN_753[31:0]; // @[programmableCache.scala 138:33 programmableCache.scala 417:31]
  wire  _T_451 = actionReg_3_io_deq_bits_action_actionType == 4'h3; // @[programmableCache.scala 373:73]
  wire  isStateAction_3 = _T_451 & actionReg_3_io_deq_valid; // @[programmableCache.scala 373:82]
  wire [1:0] tbeAction_3 = actionReg_3_io_deq_bits_action_signals[1:0]; // @[Gem5CacheLogic.scala 115:54]
  wire  _T_445 = actionReg_3_io_deq_bits_action_actionType == 4'h1; // @[programmableCache.scala 370:73]
  wire  isTBEAction_3 = _T_445 & actionReg_3_io_deq_valid; // @[programmableCache.scala 370:82]
  wire  maskField_4 = actionReg_4_io_deq_bits_action_signals[2]; // @[Gem5CacheLogic.scala 114:54]
  wire  _T_209 = ~maskField_4; // @[programmableCache.scala 303:84]
  wire [63:0] _GEN_931 = compUnit_4_io_reg_file_0; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_932 = 2'h1 == actionReg_4_io_deq_bits_action_signals[4:3] ? compUnit_4_io_reg_file_1 : _GEN_931; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_933 = 2'h2 == actionReg_4_io_deq_bits_action_signals[4:3] ? compUnit_4_io_reg_file_2 : _GEN_932; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_934 = 2'h3 == actionReg_4_io_deq_bits_action_signals[4:3] ? compUnit_4_io_reg_file_3 : _GEN_933; // @[programmableCache.scala 417:31]
  wire [31:0] tbeFieldUpdateSrc_4 = _GEN_934[31:0]; // @[programmableCache.scala 138:33 programmableCache.scala 417:31]
  wire  _T_508 = actionReg_4_io_deq_bits_action_actionType == 4'h3; // @[programmableCache.scala 373:73]
  wire  isStateAction_4 = _T_508 & actionReg_4_io_deq_valid; // @[programmableCache.scala 373:82]
  wire [1:0] tbeAction_4 = actionReg_4_io_deq_bits_action_signals[1:0]; // @[Gem5CacheLogic.scala 115:54]
  wire  _T_502 = actionReg_4_io_deq_bits_action_actionType == 4'h1; // @[programmableCache.scala 370:73]
  wire  isTBEAction_4 = _T_502 & actionReg_4_io_deq_valid; // @[programmableCache.scala 370:82]
  wire  maskField_5 = actionReg_5_io_deq_bits_action_signals[2]; // @[Gem5CacheLogic.scala 114:54]
  wire  _T_215 = ~maskField_5; // @[programmableCache.scala 303:84]
  wire [63:0] _GEN_1112 = compUnit_5_io_reg_file_0; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_1113 = 2'h1 == actionReg_5_io_deq_bits_action_signals[4:3] ? compUnit_5_io_reg_file_1 : _GEN_1112; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_1114 = 2'h2 == actionReg_5_io_deq_bits_action_signals[4:3] ? compUnit_5_io_reg_file_2 : _GEN_1113; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_1115 = 2'h3 == actionReg_5_io_deq_bits_action_signals[4:3] ? compUnit_5_io_reg_file_3 : _GEN_1114; // @[programmableCache.scala 417:31]
  wire [31:0] tbeFieldUpdateSrc_5 = _GEN_1115[31:0]; // @[programmableCache.scala 138:33 programmableCache.scala 417:31]
  wire  _T_565 = actionReg_5_io_deq_bits_action_actionType == 4'h3; // @[programmableCache.scala 373:73]
  wire  isStateAction_5 = _T_565 & actionReg_5_io_deq_valid; // @[programmableCache.scala 373:82]
  wire [1:0] tbeAction_5 = actionReg_5_io_deq_bits_action_signals[1:0]; // @[Gem5CacheLogic.scala 115:54]
  wire  _T_559 = actionReg_5_io_deq_bits_action_actionType == 4'h1; // @[programmableCache.scala 370:73]
  wire  isTBEAction_5 = _T_559 & actionReg_5_io_deq_valid; // @[programmableCache.scala 370:82]
  wire  maskField_6 = actionReg_6_io_deq_bits_action_signals[2]; // @[Gem5CacheLogic.scala 114:54]
  wire  _T_221 = ~maskField_6; // @[programmableCache.scala 303:84]
  wire [63:0] _GEN_1293 = compUnit_6_io_reg_file_0; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_1294 = 2'h1 == actionReg_6_io_deq_bits_action_signals[4:3] ? compUnit_6_io_reg_file_1 : _GEN_1293; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_1295 = 2'h2 == actionReg_6_io_deq_bits_action_signals[4:3] ? compUnit_6_io_reg_file_2 : _GEN_1294; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_1296 = 2'h3 == actionReg_6_io_deq_bits_action_signals[4:3] ? compUnit_6_io_reg_file_3 : _GEN_1295; // @[programmableCache.scala 417:31]
  wire [31:0] tbeFieldUpdateSrc_6 = _GEN_1296[31:0]; // @[programmableCache.scala 138:33 programmableCache.scala 417:31]
  wire  _T_622 = actionReg_6_io_deq_bits_action_actionType == 4'h3; // @[programmableCache.scala 373:73]
  wire  isStateAction_6 = _T_622 & actionReg_6_io_deq_valid; // @[programmableCache.scala 373:82]
  wire [1:0] tbeAction_6 = actionReg_6_io_deq_bits_action_signals[1:0]; // @[Gem5CacheLogic.scala 115:54]
  wire  _T_616 = actionReg_6_io_deq_bits_action_actionType == 4'h1; // @[programmableCache.scala 370:73]
  wire  isTBEAction_6 = _T_616 & actionReg_6_io_deq_valid; // @[programmableCache.scala 370:82]
  wire  maskField_7 = actionReg_7_io_deq_bits_action_signals[2]; // @[Gem5CacheLogic.scala 114:54]
  wire  _T_227 = ~maskField_7; // @[programmableCache.scala 303:84]
  wire [63:0] _GEN_1474 = compUnit_7_io_reg_file_0; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_1475 = 2'h1 == actionReg_7_io_deq_bits_action_signals[4:3] ? compUnit_7_io_reg_file_1 : _GEN_1474; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_1476 = 2'h2 == actionReg_7_io_deq_bits_action_signals[4:3] ? compUnit_7_io_reg_file_2 : _GEN_1475; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_1477 = 2'h3 == actionReg_7_io_deq_bits_action_signals[4:3] ? compUnit_7_io_reg_file_3 : _GEN_1476; // @[programmableCache.scala 417:31]
  wire [31:0] tbeFieldUpdateSrc_7 = _GEN_1477[31:0]; // @[programmableCache.scala 138:33 programmableCache.scala 417:31]
  wire  _T_679 = actionReg_7_io_deq_bits_action_actionType == 4'h3; // @[programmableCache.scala 373:73]
  wire  isStateAction_7 = _T_679 & actionReg_7_io_deq_valid; // @[programmableCache.scala 373:82]
  wire [1:0] tbeAction_7 = actionReg_7_io_deq_bits_action_signals[1:0]; // @[Gem5CacheLogic.scala 115:54]
  wire  _T_673 = actionReg_7_io_deq_bits_action_actionType == 4'h1; // @[programmableCache.scala 370:73]
  wire  isTBEAction_7 = _T_673 & actionReg_7_io_deq_valid; // @[programmableCache.scala 370:82]
  wire [5:0] _GEN_1 = 4'h1 == routine ? 6'h0 : 6'h1; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_2 = 4'h2 == routine ? 6'h38 : _GEN_1; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_3 = 4'h3 == routine ? 6'h3a : _GEN_2; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_4 = 4'h4 == routine ? 6'h33 : _GEN_3; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_5 = 4'h5 == routine ? 6'h15 : _GEN_4; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_6 = 4'h6 == routine ? 6'h20 : _GEN_5; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_7 = 4'h7 == routine ? 6'h0 : _GEN_6; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_8 = 4'h8 == routine ? 6'h0 : _GEN_7; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_9 = 4'h9 == routine ? 6'h0 : _GEN_8; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_10 = 4'ha == routine ? 6'h0 : _GEN_9; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_11 = 4'hb == routine ? 6'h0 : _GEN_10; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_12 = 4'hc == routine ? 6'h0 : _GEN_11; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_13 = 4'hd == routine ? 6'h0 : _GEN_12; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_14 = 4'he == routine ? 6'h0 : _GEN_13; // @[programmableCache.scala 349:30]
  wire [5:0] _GEN_15 = 4'hf == routine ? 6'h0 : _GEN_14; // @[programmableCache.scala 349:30]
  wire [31:0] addrReplacer = {{31'd0}, input__io_deq_bits_inst_addr[0]}; // @[programmableCache.scala 207:28 programmableCache.scala 356:18]
  wire  _GEN_17 = addrReplacer[0] ? replStateReg_1 : replStateReg_0; // @[Replacement.scala 97:41]
  wire [1:0] _T_241 = {_GEN_17,1'h0}; // @[Cat.scala 29:58]
  wire  _T_243 = &_T_241[1]; // @[Replacement.scala 133:103]
  wire  _T_246 = ~_T_241[1]; // @[Replacement.scala 134:89]
  wire [1:0] _T_248 = {_T_246,_T_243}; // @[Cat.scala 29:58]
  wire  replacerWayWire = _T_248[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] _T_257 = 2'h1 << replacerWayWire; // @[OneHot.scala 65:12]
  wire  _T_259 = ~replacerWayWire; // @[Replacement.scala 111:25]
  wire [1:0] _T_260 = _T_241 | _T_257; // @[Replacement.scala 111:72]
  wire [1:0] _T_261 = _T_259 ? 2'h0 : _T_260; // @[Replacement.scala 111:20]
  wire  missLD = _T_156; // @[programmableCache.scala 111:22 programmableCache.scala 277:12]
  wire [2:0] tbeWay = input__io_deq_bits_tbeOut_way; // @[programmableCache.scala 294:12]
  wire  _T_263 = tbeWay == 3'h2; // @[programmableCache.scala 363:44]
  reg [2:0] wayInputCache; // @[Reg.scala 27:20]
  reg [31:0] tbeFields_0; // @[Reg.scala 27:20]
  reg [1:0] _T_270; // @[Reg.scala 27:20]
  reg [31:0] inputToPC_addr; // @[Reg.scala 27:20]
  reg [63:0] inputToPC_data; // @[Reg.scala 27:20]
  wire  _T_276 = actionReg_0_io_deq_bits_action_actionType == 4'h0; // @[programmableCache.scala 371:73]
  wire  isCacheAction_0 = _T_276 & actionReg_0_io_deq_valid; // @[programmableCache.scala 371:82]
  wire  _T_278 = actionReg_0_io_deq_bits_action_actionType == 4'h2; // @[programmableCache.scala 372:77]
  wire  _T_282 = actionReg_0_io_deq_bits_action_actionType == 4'h4; // @[programmableCache.scala 374:72]
  wire  _T_284 = actionReg_0_io_deq_bits_action_actionType >= 4'h8; // @[programmableCache.scala 375:73]
  wire [15:0] pcWire_0_pc = pc_io_read_0_out_bits_pc; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [31:0] _GEN_31 = 6'h1 == pcWire_0_pc[5:0] ? 32'h10000001 : 32'h0; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_32 = 6'h2 == pcWire_0_pc[5:0] ? 32'h34 : _GEN_31; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_33 = 6'h3 == pcWire_0_pc[5:0] ? 32'hc0000010 : _GEN_32; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_34 = 6'h4 == pcWire_0_pc[5:0] ? 32'h1000000b : _GEN_33; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_35 = 6'h5 == pcWire_0_pc[5:0] ? 32'hf0007003 : _GEN_34; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_36 = 6'h6 == pcWire_0_pc[5:0] ? 32'hf000d013 : _GEN_35; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_37 = 6'h7 == pcWire_0_pc[5:0] ? 32'h80000405 : _GEN_36; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_38 = 6'h8 == pcWire_0_pc[5:0] ? 32'hf0015013 : _GEN_37; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_39 = 6'h9 == pcWire_0_pc[5:0] ? 32'h80000405 : _GEN_38; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_40 = 6'ha == pcWire_0_pc[5:0] ? 32'h90000005 : _GEN_39; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_41 = 6'hb == pcWire_0_pc[5:0] ? 32'he07ff011 : _GEN_40; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_42 = 6'hc == pcWire_0_pc[5:0] ? 32'he06b2016 : _GEN_41; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_43 = 6'hd == pcWire_0_pc[5:0] ? 32'h10000000 : _GEN_42; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_44 = 6'he == pcWire_0_pc[5:0] ? 32'he03ff011 : _GEN_43; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_45 = 6'hf == pcWire_0_pc[5:0] ? 32'he0003404 : _GEN_44; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_46 = 6'h10 == pcWire_0_pc[5:0] ? 32'hc0000010 : _GEN_45; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_47 = 6'h11 == pcWire_0_pc[5:0] ? 32'he0800410 : _GEN_46; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_48 = 6'h12 == pcWire_0_pc[5:0] ? 32'h40000203 : _GEN_47; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_49 = 6'h13 == pcWire_0_pc[5:0] ? 32'h30000001 : _GEN_48; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_50 = 6'h14 == pcWire_0_pc[5:0] ? 32'h0 : _GEN_49; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_51 = 6'h15 == pcWire_0_pc[5:0] ? 32'hc0000037 : _GEN_50; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_52 = 6'h16 == pcWire_0_pc[5:0] ? 32'h10000000 : _GEN_51; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_53 = 6'h17 == pcWire_0_pc[5:0] ? 32'h10000002 : _GEN_52; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_54 = 6'h18 == pcWire_0_pc[5:0] ? 32'h30000000 : _GEN_53; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_55 = 6'h19 == pcWire_0_pc[5:0] ? 32'h0 : _GEN_54; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_56 = 6'h1a == pcWire_0_pc[5:0] ? 32'hc0000010 : _GEN_55; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_57 = 6'h1b == pcWire_0_pc[5:0] ? 32'he0003404 : _GEN_56; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_58 = 6'h1c == pcWire_0_pc[5:0] ? 32'ha0000010 : _GEN_57; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_59 = 6'h1d == pcWire_0_pc[5:0] ? 32'h40000203 : _GEN_58; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_60 = 6'h1e == pcWire_0_pc[5:0] ? 32'h30000002 : _GEN_59; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_61 = 6'h1f == pcWire_0_pc[5:0] ? 32'h0 : _GEN_60; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_62 = 6'h20 == pcWire_0_pc[5:0] ? 32'heffff000 : _GEN_61; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_63 = 6'h21 == pcWire_0_pc[5:0] ? 32'he0010014 : _GEN_62; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_64 = 6'h22 == pcWire_0_pc[5:0] ? 32'h80001008 : _GEN_63; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_65 = 6'h23 == pcWire_0_pc[5:0] ? 32'hc0000011 : _GEN_64; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_66 = 6'h24 == pcWire_0_pc[5:0] ? 32'h90001027 : _GEN_65; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_67 = 6'h25 == pcWire_0_pc[5:0] ? 32'h10000000 : _GEN_66; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_68 = 6'h26 == pcWire_0_pc[5:0] ? 32'h80 : _GEN_67; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_69 = 6'h27 == pcWire_0_pc[5:0] ? 32'h100 : _GEN_68; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_70 = 6'h28 == pcWire_0_pc[5:0] ? 32'he0020004 : _GEN_69; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_71 = 6'h29 == pcWire_0_pc[5:0] ? 32'hc0000011 : _GEN_70; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_72 = 6'h2a == pcWire_0_pc[5:0] ? 32'he0001820 : _GEN_71; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_73 = 6'h2b == pcWire_0_pc[5:0] ? 32'h80002436 : _GEN_72; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_74 = 6'h2c == pcWire_0_pc[5:0] ? 32'h10000000 : _GEN_73; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_75 = 6'h2d == pcWire_0_pc[5:0] ? 32'he001d403 : _GEN_74; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_76 = 6'h2e == pcWire_0_pc[5:0] ? 32'ha0000010 : _GEN_75; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_77 = 6'h2f == pcWire_0_pc[5:0] ? 32'h40000203 : _GEN_76; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_78 = 6'h30 == pcWire_0_pc[5:0] ? 32'h10000002 : _GEN_77; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_79 = 6'h31 == pcWire_0_pc[5:0] ? 32'h30000003 : _GEN_78; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_80 = 6'h32 == pcWire_0_pc[5:0] ? 32'h0 : _GEN_79; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_81 = 6'h33 == pcWire_0_pc[5:0] ? 32'h34 : _GEN_80; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_82 = 6'h34 == pcWire_0_pc[5:0] ? 32'h80 : _GEN_81; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_83 = 6'h35 == pcWire_0_pc[5:0] ? 32'h100 : _GEN_82; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_84 = 6'h36 == pcWire_0_pc[5:0] ? 32'h30000002 : _GEN_83; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_85 = 6'h37 == pcWire_0_pc[5:0] ? 32'h0 : _GEN_84; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_86 = 6'h38 == pcWire_0_pc[5:0] ? 32'h30000002 : _GEN_85; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_87 = 6'h39 == pcWire_0_pc[5:0] ? 32'h0 : _GEN_86; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_88 = 6'h3a == pcWire_0_pc[5:0] ? 32'h30000003 : _GEN_87; // @[Gem5CacheLogic.scala 110:53]
  wire  _T_299 = pc_io_read_0_out_bits_way == 2'h2; // @[programmableCache.scala 396:52]
  wire  updateWay_0 = _T_299 & cache_io_cpu_0_resp_valid; // @[programmableCache.scala 396:64]
  wire [2:0] cacheWayWire_0 = {{1'd0}, cache_io_cpu_0_resp_bits_way}; // @[programmableCache.scala 154:28 programmableCache.scala 213:25]
  wire [1:0] pcWire_0_way = pc_io_read_0_out_bits_way; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [2:0] _T_290 = updateWay_0 ? cacheWayWire_0 : {{1'd0}, pcWire_0_way}; // @[programmableCache.scala 386:45]
  wire  firstLineNextRoutine_0 = _GEN_88 == 32'h0; // @[programmableCache.scala 392:72]
  wire [15:0] _T_294 = pcWire_0_pc + 16'h1; // @[programmableCache.scala 393:81]
  wire [15:0] _T_296 = _T_294 + compUnit_0_io_pc; // @[programmableCache.scala 393:87]
  wire [2:0] _T_301 = updateWay_0 ? cacheWayWire_0 : {{1'd0}, pc_io_read_0_out_bits_way}; // @[programmableCache.scala 398:46]
  wire  _T_333 = actionReg_1_io_deq_bits_action_actionType == 4'h0; // @[programmableCache.scala 371:73]
  wire  isCacheAction_1 = _T_333 & actionReg_1_io_deq_valid; // @[programmableCache.scala 371:82]
  wire  _T_335 = actionReg_1_io_deq_bits_action_actionType == 4'h2; // @[programmableCache.scala 372:77]
  wire  _T_339 = actionReg_1_io_deq_bits_action_actionType == 4'h4; // @[programmableCache.scala 374:72]
  wire  _T_341 = actionReg_1_io_deq_bits_action_actionType >= 4'h8; // @[programmableCache.scala 375:73]
  wire [15:0] pcWire_1_pc = pc_io_read_1_out_bits_pc; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [31:0] _GEN_212 = 6'h1 == pcWire_1_pc[5:0] ? 32'h10000001 : 32'h0; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_213 = 6'h2 == pcWire_1_pc[5:0] ? 32'h34 : _GEN_212; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_214 = 6'h3 == pcWire_1_pc[5:0] ? 32'hc0000010 : _GEN_213; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_215 = 6'h4 == pcWire_1_pc[5:0] ? 32'h1000000b : _GEN_214; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_216 = 6'h5 == pcWire_1_pc[5:0] ? 32'hf0007003 : _GEN_215; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_217 = 6'h6 == pcWire_1_pc[5:0] ? 32'hf000d013 : _GEN_216; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_218 = 6'h7 == pcWire_1_pc[5:0] ? 32'h80000405 : _GEN_217; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_219 = 6'h8 == pcWire_1_pc[5:0] ? 32'hf0015013 : _GEN_218; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_220 = 6'h9 == pcWire_1_pc[5:0] ? 32'h80000405 : _GEN_219; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_221 = 6'ha == pcWire_1_pc[5:0] ? 32'h90000005 : _GEN_220; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_222 = 6'hb == pcWire_1_pc[5:0] ? 32'he07ff011 : _GEN_221; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_223 = 6'hc == pcWire_1_pc[5:0] ? 32'he06b2016 : _GEN_222; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_224 = 6'hd == pcWire_1_pc[5:0] ? 32'h10000000 : _GEN_223; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_225 = 6'he == pcWire_1_pc[5:0] ? 32'he03ff011 : _GEN_224; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_226 = 6'hf == pcWire_1_pc[5:0] ? 32'he0003404 : _GEN_225; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_227 = 6'h10 == pcWire_1_pc[5:0] ? 32'hc0000010 : _GEN_226; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_228 = 6'h11 == pcWire_1_pc[5:0] ? 32'he0800410 : _GEN_227; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_229 = 6'h12 == pcWire_1_pc[5:0] ? 32'h40000203 : _GEN_228; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_230 = 6'h13 == pcWire_1_pc[5:0] ? 32'h30000001 : _GEN_229; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_231 = 6'h14 == pcWire_1_pc[5:0] ? 32'h0 : _GEN_230; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_232 = 6'h15 == pcWire_1_pc[5:0] ? 32'hc0000037 : _GEN_231; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_233 = 6'h16 == pcWire_1_pc[5:0] ? 32'h10000000 : _GEN_232; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_234 = 6'h17 == pcWire_1_pc[5:0] ? 32'h10000002 : _GEN_233; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_235 = 6'h18 == pcWire_1_pc[5:0] ? 32'h30000000 : _GEN_234; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_236 = 6'h19 == pcWire_1_pc[5:0] ? 32'h0 : _GEN_235; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_237 = 6'h1a == pcWire_1_pc[5:0] ? 32'hc0000010 : _GEN_236; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_238 = 6'h1b == pcWire_1_pc[5:0] ? 32'he0003404 : _GEN_237; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_239 = 6'h1c == pcWire_1_pc[5:0] ? 32'ha0000010 : _GEN_238; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_240 = 6'h1d == pcWire_1_pc[5:0] ? 32'h40000203 : _GEN_239; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_241 = 6'h1e == pcWire_1_pc[5:0] ? 32'h30000002 : _GEN_240; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_242 = 6'h1f == pcWire_1_pc[5:0] ? 32'h0 : _GEN_241; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_243 = 6'h20 == pcWire_1_pc[5:0] ? 32'heffff000 : _GEN_242; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_244 = 6'h21 == pcWire_1_pc[5:0] ? 32'he0010014 : _GEN_243; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_245 = 6'h22 == pcWire_1_pc[5:0] ? 32'h80001008 : _GEN_244; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_246 = 6'h23 == pcWire_1_pc[5:0] ? 32'hc0000011 : _GEN_245; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_247 = 6'h24 == pcWire_1_pc[5:0] ? 32'h90001027 : _GEN_246; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_248 = 6'h25 == pcWire_1_pc[5:0] ? 32'h10000000 : _GEN_247; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_249 = 6'h26 == pcWire_1_pc[5:0] ? 32'h80 : _GEN_248; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_250 = 6'h27 == pcWire_1_pc[5:0] ? 32'h100 : _GEN_249; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_251 = 6'h28 == pcWire_1_pc[5:0] ? 32'he0020004 : _GEN_250; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_252 = 6'h29 == pcWire_1_pc[5:0] ? 32'hc0000011 : _GEN_251; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_253 = 6'h2a == pcWire_1_pc[5:0] ? 32'he0001820 : _GEN_252; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_254 = 6'h2b == pcWire_1_pc[5:0] ? 32'h80002436 : _GEN_253; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_255 = 6'h2c == pcWire_1_pc[5:0] ? 32'h10000000 : _GEN_254; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_256 = 6'h2d == pcWire_1_pc[5:0] ? 32'he001d403 : _GEN_255; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_257 = 6'h2e == pcWire_1_pc[5:0] ? 32'ha0000010 : _GEN_256; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_258 = 6'h2f == pcWire_1_pc[5:0] ? 32'h40000203 : _GEN_257; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_259 = 6'h30 == pcWire_1_pc[5:0] ? 32'h10000002 : _GEN_258; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_260 = 6'h31 == pcWire_1_pc[5:0] ? 32'h30000003 : _GEN_259; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_261 = 6'h32 == pcWire_1_pc[5:0] ? 32'h0 : _GEN_260; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_262 = 6'h33 == pcWire_1_pc[5:0] ? 32'h34 : _GEN_261; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_263 = 6'h34 == pcWire_1_pc[5:0] ? 32'h80 : _GEN_262; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_264 = 6'h35 == pcWire_1_pc[5:0] ? 32'h100 : _GEN_263; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_265 = 6'h36 == pcWire_1_pc[5:0] ? 32'h30000002 : _GEN_264; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_266 = 6'h37 == pcWire_1_pc[5:0] ? 32'h0 : _GEN_265; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_267 = 6'h38 == pcWire_1_pc[5:0] ? 32'h30000002 : _GEN_266; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_268 = 6'h39 == pcWire_1_pc[5:0] ? 32'h0 : _GEN_267; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_269 = 6'h3a == pcWire_1_pc[5:0] ? 32'h30000003 : _GEN_268; // @[Gem5CacheLogic.scala 110:53]
  wire  _T_356 = pc_io_read_1_out_bits_way == 2'h2; // @[programmableCache.scala 396:52]
  wire  updateWay_1 = _T_356 & cache_io_cpu_1_resp_valid; // @[programmableCache.scala 396:64]
  wire [2:0] cacheWayWire_1 = {{1'd0}, cache_io_cpu_1_resp_bits_way}; // @[programmableCache.scala 154:28 programmableCache.scala 213:25]
  wire [1:0] pcWire_1_way = pc_io_read_1_out_bits_way; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [2:0] _T_347 = updateWay_1 ? cacheWayWire_1 : {{1'd0}, pcWire_1_way}; // @[programmableCache.scala 386:45]
  wire  firstLineNextRoutine_1 = _GEN_269 == 32'h0; // @[programmableCache.scala 392:72]
  wire [15:0] _T_351 = pcWire_1_pc + 16'h1; // @[programmableCache.scala 393:81]
  wire [15:0] _T_353 = _T_351 + compUnit_1_io_pc; // @[programmableCache.scala 393:87]
  wire [2:0] _T_358 = updateWay_1 ? cacheWayWire_1 : {{1'd0}, pc_io_read_1_out_bits_way}; // @[programmableCache.scala 398:46]
  wire  _T_390 = actionReg_2_io_deq_bits_action_actionType == 4'h0; // @[programmableCache.scala 371:73]
  wire  isCacheAction_2 = _T_390 & actionReg_2_io_deq_valid; // @[programmableCache.scala 371:82]
  wire  _T_392 = actionReg_2_io_deq_bits_action_actionType == 4'h2; // @[programmableCache.scala 372:77]
  wire  _T_396 = actionReg_2_io_deq_bits_action_actionType == 4'h4; // @[programmableCache.scala 374:72]
  wire  _T_398 = actionReg_2_io_deq_bits_action_actionType >= 4'h8; // @[programmableCache.scala 375:73]
  wire [15:0] pcWire_2_pc = pc_io_read_2_out_bits_pc; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [31:0] _GEN_393 = 6'h1 == pcWire_2_pc[5:0] ? 32'h10000001 : 32'h0; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_394 = 6'h2 == pcWire_2_pc[5:0] ? 32'h34 : _GEN_393; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_395 = 6'h3 == pcWire_2_pc[5:0] ? 32'hc0000010 : _GEN_394; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_396 = 6'h4 == pcWire_2_pc[5:0] ? 32'h1000000b : _GEN_395; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_397 = 6'h5 == pcWire_2_pc[5:0] ? 32'hf0007003 : _GEN_396; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_398 = 6'h6 == pcWire_2_pc[5:0] ? 32'hf000d013 : _GEN_397; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_399 = 6'h7 == pcWire_2_pc[5:0] ? 32'h80000405 : _GEN_398; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_400 = 6'h8 == pcWire_2_pc[5:0] ? 32'hf0015013 : _GEN_399; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_401 = 6'h9 == pcWire_2_pc[5:0] ? 32'h80000405 : _GEN_400; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_402 = 6'ha == pcWire_2_pc[5:0] ? 32'h90000005 : _GEN_401; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_403 = 6'hb == pcWire_2_pc[5:0] ? 32'he07ff011 : _GEN_402; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_404 = 6'hc == pcWire_2_pc[5:0] ? 32'he06b2016 : _GEN_403; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_405 = 6'hd == pcWire_2_pc[5:0] ? 32'h10000000 : _GEN_404; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_406 = 6'he == pcWire_2_pc[5:0] ? 32'he03ff011 : _GEN_405; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_407 = 6'hf == pcWire_2_pc[5:0] ? 32'he0003404 : _GEN_406; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_408 = 6'h10 == pcWire_2_pc[5:0] ? 32'hc0000010 : _GEN_407; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_409 = 6'h11 == pcWire_2_pc[5:0] ? 32'he0800410 : _GEN_408; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_410 = 6'h12 == pcWire_2_pc[5:0] ? 32'h40000203 : _GEN_409; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_411 = 6'h13 == pcWire_2_pc[5:0] ? 32'h30000001 : _GEN_410; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_412 = 6'h14 == pcWire_2_pc[5:0] ? 32'h0 : _GEN_411; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_413 = 6'h15 == pcWire_2_pc[5:0] ? 32'hc0000037 : _GEN_412; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_414 = 6'h16 == pcWire_2_pc[5:0] ? 32'h10000000 : _GEN_413; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_415 = 6'h17 == pcWire_2_pc[5:0] ? 32'h10000002 : _GEN_414; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_416 = 6'h18 == pcWire_2_pc[5:0] ? 32'h30000000 : _GEN_415; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_417 = 6'h19 == pcWire_2_pc[5:0] ? 32'h0 : _GEN_416; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_418 = 6'h1a == pcWire_2_pc[5:0] ? 32'hc0000010 : _GEN_417; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_419 = 6'h1b == pcWire_2_pc[5:0] ? 32'he0003404 : _GEN_418; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_420 = 6'h1c == pcWire_2_pc[5:0] ? 32'ha0000010 : _GEN_419; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_421 = 6'h1d == pcWire_2_pc[5:0] ? 32'h40000203 : _GEN_420; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_422 = 6'h1e == pcWire_2_pc[5:0] ? 32'h30000002 : _GEN_421; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_423 = 6'h1f == pcWire_2_pc[5:0] ? 32'h0 : _GEN_422; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_424 = 6'h20 == pcWire_2_pc[5:0] ? 32'heffff000 : _GEN_423; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_425 = 6'h21 == pcWire_2_pc[5:0] ? 32'he0010014 : _GEN_424; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_426 = 6'h22 == pcWire_2_pc[5:0] ? 32'h80001008 : _GEN_425; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_427 = 6'h23 == pcWire_2_pc[5:0] ? 32'hc0000011 : _GEN_426; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_428 = 6'h24 == pcWire_2_pc[5:0] ? 32'h90001027 : _GEN_427; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_429 = 6'h25 == pcWire_2_pc[5:0] ? 32'h10000000 : _GEN_428; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_430 = 6'h26 == pcWire_2_pc[5:0] ? 32'h80 : _GEN_429; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_431 = 6'h27 == pcWire_2_pc[5:0] ? 32'h100 : _GEN_430; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_432 = 6'h28 == pcWire_2_pc[5:0] ? 32'he0020004 : _GEN_431; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_433 = 6'h29 == pcWire_2_pc[5:0] ? 32'hc0000011 : _GEN_432; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_434 = 6'h2a == pcWire_2_pc[5:0] ? 32'he0001820 : _GEN_433; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_435 = 6'h2b == pcWire_2_pc[5:0] ? 32'h80002436 : _GEN_434; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_436 = 6'h2c == pcWire_2_pc[5:0] ? 32'h10000000 : _GEN_435; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_437 = 6'h2d == pcWire_2_pc[5:0] ? 32'he001d403 : _GEN_436; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_438 = 6'h2e == pcWire_2_pc[5:0] ? 32'ha0000010 : _GEN_437; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_439 = 6'h2f == pcWire_2_pc[5:0] ? 32'h40000203 : _GEN_438; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_440 = 6'h30 == pcWire_2_pc[5:0] ? 32'h10000002 : _GEN_439; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_441 = 6'h31 == pcWire_2_pc[5:0] ? 32'h30000003 : _GEN_440; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_442 = 6'h32 == pcWire_2_pc[5:0] ? 32'h0 : _GEN_441; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_443 = 6'h33 == pcWire_2_pc[5:0] ? 32'h34 : _GEN_442; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_444 = 6'h34 == pcWire_2_pc[5:0] ? 32'h80 : _GEN_443; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_445 = 6'h35 == pcWire_2_pc[5:0] ? 32'h100 : _GEN_444; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_446 = 6'h36 == pcWire_2_pc[5:0] ? 32'h30000002 : _GEN_445; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_447 = 6'h37 == pcWire_2_pc[5:0] ? 32'h0 : _GEN_446; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_448 = 6'h38 == pcWire_2_pc[5:0] ? 32'h30000002 : _GEN_447; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_449 = 6'h39 == pcWire_2_pc[5:0] ? 32'h0 : _GEN_448; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_450 = 6'h3a == pcWire_2_pc[5:0] ? 32'h30000003 : _GEN_449; // @[Gem5CacheLogic.scala 110:53]
  wire  _T_413 = pc_io_read_2_out_bits_way == 2'h2; // @[programmableCache.scala 396:52]
  wire  updateWay_2 = _T_413 & cache_io_cpu_2_resp_valid; // @[programmableCache.scala 396:64]
  wire [2:0] cacheWayWire_2 = {{1'd0}, cache_io_cpu_2_resp_bits_way}; // @[programmableCache.scala 154:28 programmableCache.scala 213:25]
  wire [1:0] pcWire_2_way = pc_io_read_2_out_bits_way; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [2:0] _T_404 = updateWay_2 ? cacheWayWire_2 : {{1'd0}, pcWire_2_way}; // @[programmableCache.scala 386:45]
  wire  firstLineNextRoutine_2 = _GEN_450 == 32'h0; // @[programmableCache.scala 392:72]
  wire [15:0] _T_408 = pcWire_2_pc + 16'h1; // @[programmableCache.scala 393:81]
  wire [15:0] _T_410 = _T_408 + compUnit_2_io_pc; // @[programmableCache.scala 393:87]
  wire [2:0] _T_415 = updateWay_2 ? cacheWayWire_2 : {{1'd0}, pc_io_read_2_out_bits_way}; // @[programmableCache.scala 398:46]
  wire  _T_447 = actionReg_3_io_deq_bits_action_actionType == 4'h0; // @[programmableCache.scala 371:73]
  wire  isCacheAction_3 = _T_447 & actionReg_3_io_deq_valid; // @[programmableCache.scala 371:82]
  wire  _T_449 = actionReg_3_io_deq_bits_action_actionType == 4'h2; // @[programmableCache.scala 372:77]
  wire  _T_453 = actionReg_3_io_deq_bits_action_actionType == 4'h4; // @[programmableCache.scala 374:72]
  wire  _T_455 = actionReg_3_io_deq_bits_action_actionType >= 4'h8; // @[programmableCache.scala 375:73]
  wire [15:0] pcWire_3_pc = pc_io_read_3_out_bits_pc; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [31:0] _GEN_574 = 6'h1 == pcWire_3_pc[5:0] ? 32'h10000001 : 32'h0; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_575 = 6'h2 == pcWire_3_pc[5:0] ? 32'h34 : _GEN_574; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_576 = 6'h3 == pcWire_3_pc[5:0] ? 32'hc0000010 : _GEN_575; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_577 = 6'h4 == pcWire_3_pc[5:0] ? 32'h1000000b : _GEN_576; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_578 = 6'h5 == pcWire_3_pc[5:0] ? 32'hf0007003 : _GEN_577; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_579 = 6'h6 == pcWire_3_pc[5:0] ? 32'hf000d013 : _GEN_578; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_580 = 6'h7 == pcWire_3_pc[5:0] ? 32'h80000405 : _GEN_579; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_581 = 6'h8 == pcWire_3_pc[5:0] ? 32'hf0015013 : _GEN_580; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_582 = 6'h9 == pcWire_3_pc[5:0] ? 32'h80000405 : _GEN_581; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_583 = 6'ha == pcWire_3_pc[5:0] ? 32'h90000005 : _GEN_582; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_584 = 6'hb == pcWire_3_pc[5:0] ? 32'he07ff011 : _GEN_583; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_585 = 6'hc == pcWire_3_pc[5:0] ? 32'he06b2016 : _GEN_584; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_586 = 6'hd == pcWire_3_pc[5:0] ? 32'h10000000 : _GEN_585; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_587 = 6'he == pcWire_3_pc[5:0] ? 32'he03ff011 : _GEN_586; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_588 = 6'hf == pcWire_3_pc[5:0] ? 32'he0003404 : _GEN_587; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_589 = 6'h10 == pcWire_3_pc[5:0] ? 32'hc0000010 : _GEN_588; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_590 = 6'h11 == pcWire_3_pc[5:0] ? 32'he0800410 : _GEN_589; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_591 = 6'h12 == pcWire_3_pc[5:0] ? 32'h40000203 : _GEN_590; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_592 = 6'h13 == pcWire_3_pc[5:0] ? 32'h30000001 : _GEN_591; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_593 = 6'h14 == pcWire_3_pc[5:0] ? 32'h0 : _GEN_592; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_594 = 6'h15 == pcWire_3_pc[5:0] ? 32'hc0000037 : _GEN_593; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_595 = 6'h16 == pcWire_3_pc[5:0] ? 32'h10000000 : _GEN_594; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_596 = 6'h17 == pcWire_3_pc[5:0] ? 32'h10000002 : _GEN_595; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_597 = 6'h18 == pcWire_3_pc[5:0] ? 32'h30000000 : _GEN_596; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_598 = 6'h19 == pcWire_3_pc[5:0] ? 32'h0 : _GEN_597; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_599 = 6'h1a == pcWire_3_pc[5:0] ? 32'hc0000010 : _GEN_598; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_600 = 6'h1b == pcWire_3_pc[5:0] ? 32'he0003404 : _GEN_599; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_601 = 6'h1c == pcWire_3_pc[5:0] ? 32'ha0000010 : _GEN_600; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_602 = 6'h1d == pcWire_3_pc[5:0] ? 32'h40000203 : _GEN_601; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_603 = 6'h1e == pcWire_3_pc[5:0] ? 32'h30000002 : _GEN_602; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_604 = 6'h1f == pcWire_3_pc[5:0] ? 32'h0 : _GEN_603; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_605 = 6'h20 == pcWire_3_pc[5:0] ? 32'heffff000 : _GEN_604; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_606 = 6'h21 == pcWire_3_pc[5:0] ? 32'he0010014 : _GEN_605; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_607 = 6'h22 == pcWire_3_pc[5:0] ? 32'h80001008 : _GEN_606; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_608 = 6'h23 == pcWire_3_pc[5:0] ? 32'hc0000011 : _GEN_607; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_609 = 6'h24 == pcWire_3_pc[5:0] ? 32'h90001027 : _GEN_608; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_610 = 6'h25 == pcWire_3_pc[5:0] ? 32'h10000000 : _GEN_609; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_611 = 6'h26 == pcWire_3_pc[5:0] ? 32'h80 : _GEN_610; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_612 = 6'h27 == pcWire_3_pc[5:0] ? 32'h100 : _GEN_611; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_613 = 6'h28 == pcWire_3_pc[5:0] ? 32'he0020004 : _GEN_612; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_614 = 6'h29 == pcWire_3_pc[5:0] ? 32'hc0000011 : _GEN_613; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_615 = 6'h2a == pcWire_3_pc[5:0] ? 32'he0001820 : _GEN_614; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_616 = 6'h2b == pcWire_3_pc[5:0] ? 32'h80002436 : _GEN_615; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_617 = 6'h2c == pcWire_3_pc[5:0] ? 32'h10000000 : _GEN_616; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_618 = 6'h2d == pcWire_3_pc[5:0] ? 32'he001d403 : _GEN_617; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_619 = 6'h2e == pcWire_3_pc[5:0] ? 32'ha0000010 : _GEN_618; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_620 = 6'h2f == pcWire_3_pc[5:0] ? 32'h40000203 : _GEN_619; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_621 = 6'h30 == pcWire_3_pc[5:0] ? 32'h10000002 : _GEN_620; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_622 = 6'h31 == pcWire_3_pc[5:0] ? 32'h30000003 : _GEN_621; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_623 = 6'h32 == pcWire_3_pc[5:0] ? 32'h0 : _GEN_622; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_624 = 6'h33 == pcWire_3_pc[5:0] ? 32'h34 : _GEN_623; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_625 = 6'h34 == pcWire_3_pc[5:0] ? 32'h80 : _GEN_624; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_626 = 6'h35 == pcWire_3_pc[5:0] ? 32'h100 : _GEN_625; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_627 = 6'h36 == pcWire_3_pc[5:0] ? 32'h30000002 : _GEN_626; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_628 = 6'h37 == pcWire_3_pc[5:0] ? 32'h0 : _GEN_627; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_629 = 6'h38 == pcWire_3_pc[5:0] ? 32'h30000002 : _GEN_628; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_630 = 6'h39 == pcWire_3_pc[5:0] ? 32'h0 : _GEN_629; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_631 = 6'h3a == pcWire_3_pc[5:0] ? 32'h30000003 : _GEN_630; // @[Gem5CacheLogic.scala 110:53]
  wire  _T_470 = pc_io_read_3_out_bits_way == 2'h2; // @[programmableCache.scala 396:52]
  wire  updateWay_3 = _T_470 & cache_io_cpu_3_resp_valid; // @[programmableCache.scala 396:64]
  wire [2:0] cacheWayWire_3 = {{1'd0}, cache_io_cpu_3_resp_bits_way}; // @[programmableCache.scala 154:28 programmableCache.scala 213:25]
  wire [1:0] pcWire_3_way = pc_io_read_3_out_bits_way; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [2:0] _T_461 = updateWay_3 ? cacheWayWire_3 : {{1'd0}, pcWire_3_way}; // @[programmableCache.scala 386:45]
  wire  firstLineNextRoutine_3 = _GEN_631 == 32'h0; // @[programmableCache.scala 392:72]
  wire [15:0] _T_465 = pcWire_3_pc + 16'h1; // @[programmableCache.scala 393:81]
  wire [15:0] _T_467 = _T_465 + compUnit_3_io_pc; // @[programmableCache.scala 393:87]
  wire [2:0] _T_472 = updateWay_3 ? cacheWayWire_3 : {{1'd0}, pc_io_read_3_out_bits_way}; // @[programmableCache.scala 398:46]
  wire  _T_504 = actionReg_4_io_deq_bits_action_actionType == 4'h0; // @[programmableCache.scala 371:73]
  wire  isCacheAction_4 = _T_504 & actionReg_4_io_deq_valid; // @[programmableCache.scala 371:82]
  wire  _T_506 = actionReg_4_io_deq_bits_action_actionType == 4'h2; // @[programmableCache.scala 372:77]
  wire  _T_510 = actionReg_4_io_deq_bits_action_actionType == 4'h4; // @[programmableCache.scala 374:72]
  wire  _T_512 = actionReg_4_io_deq_bits_action_actionType >= 4'h8; // @[programmableCache.scala 375:73]
  wire [15:0] pcWire_4_pc = pc_io_read_4_out_bits_pc; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [31:0] _GEN_755 = 6'h1 == pcWire_4_pc[5:0] ? 32'h10000001 : 32'h0; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_756 = 6'h2 == pcWire_4_pc[5:0] ? 32'h34 : _GEN_755; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_757 = 6'h3 == pcWire_4_pc[5:0] ? 32'hc0000010 : _GEN_756; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_758 = 6'h4 == pcWire_4_pc[5:0] ? 32'h1000000b : _GEN_757; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_759 = 6'h5 == pcWire_4_pc[5:0] ? 32'hf0007003 : _GEN_758; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_760 = 6'h6 == pcWire_4_pc[5:0] ? 32'hf000d013 : _GEN_759; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_761 = 6'h7 == pcWire_4_pc[5:0] ? 32'h80000405 : _GEN_760; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_762 = 6'h8 == pcWire_4_pc[5:0] ? 32'hf0015013 : _GEN_761; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_763 = 6'h9 == pcWire_4_pc[5:0] ? 32'h80000405 : _GEN_762; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_764 = 6'ha == pcWire_4_pc[5:0] ? 32'h90000005 : _GEN_763; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_765 = 6'hb == pcWire_4_pc[5:0] ? 32'he07ff011 : _GEN_764; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_766 = 6'hc == pcWire_4_pc[5:0] ? 32'he06b2016 : _GEN_765; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_767 = 6'hd == pcWire_4_pc[5:0] ? 32'h10000000 : _GEN_766; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_768 = 6'he == pcWire_4_pc[5:0] ? 32'he03ff011 : _GEN_767; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_769 = 6'hf == pcWire_4_pc[5:0] ? 32'he0003404 : _GEN_768; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_770 = 6'h10 == pcWire_4_pc[5:0] ? 32'hc0000010 : _GEN_769; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_771 = 6'h11 == pcWire_4_pc[5:0] ? 32'he0800410 : _GEN_770; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_772 = 6'h12 == pcWire_4_pc[5:0] ? 32'h40000203 : _GEN_771; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_773 = 6'h13 == pcWire_4_pc[5:0] ? 32'h30000001 : _GEN_772; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_774 = 6'h14 == pcWire_4_pc[5:0] ? 32'h0 : _GEN_773; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_775 = 6'h15 == pcWire_4_pc[5:0] ? 32'hc0000037 : _GEN_774; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_776 = 6'h16 == pcWire_4_pc[5:0] ? 32'h10000000 : _GEN_775; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_777 = 6'h17 == pcWire_4_pc[5:0] ? 32'h10000002 : _GEN_776; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_778 = 6'h18 == pcWire_4_pc[5:0] ? 32'h30000000 : _GEN_777; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_779 = 6'h19 == pcWire_4_pc[5:0] ? 32'h0 : _GEN_778; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_780 = 6'h1a == pcWire_4_pc[5:0] ? 32'hc0000010 : _GEN_779; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_781 = 6'h1b == pcWire_4_pc[5:0] ? 32'he0003404 : _GEN_780; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_782 = 6'h1c == pcWire_4_pc[5:0] ? 32'ha0000010 : _GEN_781; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_783 = 6'h1d == pcWire_4_pc[5:0] ? 32'h40000203 : _GEN_782; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_784 = 6'h1e == pcWire_4_pc[5:0] ? 32'h30000002 : _GEN_783; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_785 = 6'h1f == pcWire_4_pc[5:0] ? 32'h0 : _GEN_784; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_786 = 6'h20 == pcWire_4_pc[5:0] ? 32'heffff000 : _GEN_785; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_787 = 6'h21 == pcWire_4_pc[5:0] ? 32'he0010014 : _GEN_786; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_788 = 6'h22 == pcWire_4_pc[5:0] ? 32'h80001008 : _GEN_787; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_789 = 6'h23 == pcWire_4_pc[5:0] ? 32'hc0000011 : _GEN_788; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_790 = 6'h24 == pcWire_4_pc[5:0] ? 32'h90001027 : _GEN_789; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_791 = 6'h25 == pcWire_4_pc[5:0] ? 32'h10000000 : _GEN_790; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_792 = 6'h26 == pcWire_4_pc[5:0] ? 32'h80 : _GEN_791; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_793 = 6'h27 == pcWire_4_pc[5:0] ? 32'h100 : _GEN_792; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_794 = 6'h28 == pcWire_4_pc[5:0] ? 32'he0020004 : _GEN_793; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_795 = 6'h29 == pcWire_4_pc[5:0] ? 32'hc0000011 : _GEN_794; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_796 = 6'h2a == pcWire_4_pc[5:0] ? 32'he0001820 : _GEN_795; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_797 = 6'h2b == pcWire_4_pc[5:0] ? 32'h80002436 : _GEN_796; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_798 = 6'h2c == pcWire_4_pc[5:0] ? 32'h10000000 : _GEN_797; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_799 = 6'h2d == pcWire_4_pc[5:0] ? 32'he001d403 : _GEN_798; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_800 = 6'h2e == pcWire_4_pc[5:0] ? 32'ha0000010 : _GEN_799; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_801 = 6'h2f == pcWire_4_pc[5:0] ? 32'h40000203 : _GEN_800; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_802 = 6'h30 == pcWire_4_pc[5:0] ? 32'h10000002 : _GEN_801; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_803 = 6'h31 == pcWire_4_pc[5:0] ? 32'h30000003 : _GEN_802; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_804 = 6'h32 == pcWire_4_pc[5:0] ? 32'h0 : _GEN_803; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_805 = 6'h33 == pcWire_4_pc[5:0] ? 32'h34 : _GEN_804; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_806 = 6'h34 == pcWire_4_pc[5:0] ? 32'h80 : _GEN_805; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_807 = 6'h35 == pcWire_4_pc[5:0] ? 32'h100 : _GEN_806; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_808 = 6'h36 == pcWire_4_pc[5:0] ? 32'h30000002 : _GEN_807; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_809 = 6'h37 == pcWire_4_pc[5:0] ? 32'h0 : _GEN_808; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_810 = 6'h38 == pcWire_4_pc[5:0] ? 32'h30000002 : _GEN_809; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_811 = 6'h39 == pcWire_4_pc[5:0] ? 32'h0 : _GEN_810; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_812 = 6'h3a == pcWire_4_pc[5:0] ? 32'h30000003 : _GEN_811; // @[Gem5CacheLogic.scala 110:53]
  wire  _T_527 = pc_io_read_4_out_bits_way == 2'h2; // @[programmableCache.scala 396:52]
  wire  updateWay_4 = _T_527 & cache_io_cpu_4_resp_valid; // @[programmableCache.scala 396:64]
  wire [2:0] cacheWayWire_4 = {{1'd0}, cache_io_cpu_4_resp_bits_way}; // @[programmableCache.scala 154:28 programmableCache.scala 213:25]
  wire [1:0] pcWire_4_way = pc_io_read_4_out_bits_way; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [2:0] _T_518 = updateWay_4 ? cacheWayWire_4 : {{1'd0}, pcWire_4_way}; // @[programmableCache.scala 386:45]
  wire  firstLineNextRoutine_4 = _GEN_812 == 32'h0; // @[programmableCache.scala 392:72]
  wire [15:0] _T_522 = pcWire_4_pc + 16'h1; // @[programmableCache.scala 393:81]
  wire [15:0] _T_524 = _T_522 + compUnit_4_io_pc; // @[programmableCache.scala 393:87]
  wire [2:0] _T_529 = updateWay_4 ? cacheWayWire_4 : {{1'd0}, pc_io_read_4_out_bits_way}; // @[programmableCache.scala 398:46]
  wire  _T_561 = actionReg_5_io_deq_bits_action_actionType == 4'h0; // @[programmableCache.scala 371:73]
  wire  isCacheAction_5 = _T_561 & actionReg_5_io_deq_valid; // @[programmableCache.scala 371:82]
  wire  _T_563 = actionReg_5_io_deq_bits_action_actionType == 4'h2; // @[programmableCache.scala 372:77]
  wire  _T_567 = actionReg_5_io_deq_bits_action_actionType == 4'h4; // @[programmableCache.scala 374:72]
  wire  _T_569 = actionReg_5_io_deq_bits_action_actionType >= 4'h8; // @[programmableCache.scala 375:73]
  wire [15:0] pcWire_5_pc = pc_io_read_5_out_bits_pc; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [31:0] _GEN_936 = 6'h1 == pcWire_5_pc[5:0] ? 32'h10000001 : 32'h0; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_937 = 6'h2 == pcWire_5_pc[5:0] ? 32'h34 : _GEN_936; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_938 = 6'h3 == pcWire_5_pc[5:0] ? 32'hc0000010 : _GEN_937; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_939 = 6'h4 == pcWire_5_pc[5:0] ? 32'h1000000b : _GEN_938; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_940 = 6'h5 == pcWire_5_pc[5:0] ? 32'hf0007003 : _GEN_939; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_941 = 6'h6 == pcWire_5_pc[5:0] ? 32'hf000d013 : _GEN_940; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_942 = 6'h7 == pcWire_5_pc[5:0] ? 32'h80000405 : _GEN_941; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_943 = 6'h8 == pcWire_5_pc[5:0] ? 32'hf0015013 : _GEN_942; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_944 = 6'h9 == pcWire_5_pc[5:0] ? 32'h80000405 : _GEN_943; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_945 = 6'ha == pcWire_5_pc[5:0] ? 32'h90000005 : _GEN_944; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_946 = 6'hb == pcWire_5_pc[5:0] ? 32'he07ff011 : _GEN_945; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_947 = 6'hc == pcWire_5_pc[5:0] ? 32'he06b2016 : _GEN_946; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_948 = 6'hd == pcWire_5_pc[5:0] ? 32'h10000000 : _GEN_947; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_949 = 6'he == pcWire_5_pc[5:0] ? 32'he03ff011 : _GEN_948; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_950 = 6'hf == pcWire_5_pc[5:0] ? 32'he0003404 : _GEN_949; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_951 = 6'h10 == pcWire_5_pc[5:0] ? 32'hc0000010 : _GEN_950; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_952 = 6'h11 == pcWire_5_pc[5:0] ? 32'he0800410 : _GEN_951; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_953 = 6'h12 == pcWire_5_pc[5:0] ? 32'h40000203 : _GEN_952; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_954 = 6'h13 == pcWire_5_pc[5:0] ? 32'h30000001 : _GEN_953; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_955 = 6'h14 == pcWire_5_pc[5:0] ? 32'h0 : _GEN_954; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_956 = 6'h15 == pcWire_5_pc[5:0] ? 32'hc0000037 : _GEN_955; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_957 = 6'h16 == pcWire_5_pc[5:0] ? 32'h10000000 : _GEN_956; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_958 = 6'h17 == pcWire_5_pc[5:0] ? 32'h10000002 : _GEN_957; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_959 = 6'h18 == pcWire_5_pc[5:0] ? 32'h30000000 : _GEN_958; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_960 = 6'h19 == pcWire_5_pc[5:0] ? 32'h0 : _GEN_959; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_961 = 6'h1a == pcWire_5_pc[5:0] ? 32'hc0000010 : _GEN_960; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_962 = 6'h1b == pcWire_5_pc[5:0] ? 32'he0003404 : _GEN_961; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_963 = 6'h1c == pcWire_5_pc[5:0] ? 32'ha0000010 : _GEN_962; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_964 = 6'h1d == pcWire_5_pc[5:0] ? 32'h40000203 : _GEN_963; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_965 = 6'h1e == pcWire_5_pc[5:0] ? 32'h30000002 : _GEN_964; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_966 = 6'h1f == pcWire_5_pc[5:0] ? 32'h0 : _GEN_965; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_967 = 6'h20 == pcWire_5_pc[5:0] ? 32'heffff000 : _GEN_966; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_968 = 6'h21 == pcWire_5_pc[5:0] ? 32'he0010014 : _GEN_967; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_969 = 6'h22 == pcWire_5_pc[5:0] ? 32'h80001008 : _GEN_968; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_970 = 6'h23 == pcWire_5_pc[5:0] ? 32'hc0000011 : _GEN_969; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_971 = 6'h24 == pcWire_5_pc[5:0] ? 32'h90001027 : _GEN_970; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_972 = 6'h25 == pcWire_5_pc[5:0] ? 32'h10000000 : _GEN_971; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_973 = 6'h26 == pcWire_5_pc[5:0] ? 32'h80 : _GEN_972; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_974 = 6'h27 == pcWire_5_pc[5:0] ? 32'h100 : _GEN_973; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_975 = 6'h28 == pcWire_5_pc[5:0] ? 32'he0020004 : _GEN_974; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_976 = 6'h29 == pcWire_5_pc[5:0] ? 32'hc0000011 : _GEN_975; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_977 = 6'h2a == pcWire_5_pc[5:0] ? 32'he0001820 : _GEN_976; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_978 = 6'h2b == pcWire_5_pc[5:0] ? 32'h80002436 : _GEN_977; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_979 = 6'h2c == pcWire_5_pc[5:0] ? 32'h10000000 : _GEN_978; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_980 = 6'h2d == pcWire_5_pc[5:0] ? 32'he001d403 : _GEN_979; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_981 = 6'h2e == pcWire_5_pc[5:0] ? 32'ha0000010 : _GEN_980; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_982 = 6'h2f == pcWire_5_pc[5:0] ? 32'h40000203 : _GEN_981; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_983 = 6'h30 == pcWire_5_pc[5:0] ? 32'h10000002 : _GEN_982; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_984 = 6'h31 == pcWire_5_pc[5:0] ? 32'h30000003 : _GEN_983; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_985 = 6'h32 == pcWire_5_pc[5:0] ? 32'h0 : _GEN_984; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_986 = 6'h33 == pcWire_5_pc[5:0] ? 32'h34 : _GEN_985; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_987 = 6'h34 == pcWire_5_pc[5:0] ? 32'h80 : _GEN_986; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_988 = 6'h35 == pcWire_5_pc[5:0] ? 32'h100 : _GEN_987; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_989 = 6'h36 == pcWire_5_pc[5:0] ? 32'h30000002 : _GEN_988; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_990 = 6'h37 == pcWire_5_pc[5:0] ? 32'h0 : _GEN_989; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_991 = 6'h38 == pcWire_5_pc[5:0] ? 32'h30000002 : _GEN_990; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_992 = 6'h39 == pcWire_5_pc[5:0] ? 32'h0 : _GEN_991; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_993 = 6'h3a == pcWire_5_pc[5:0] ? 32'h30000003 : _GEN_992; // @[Gem5CacheLogic.scala 110:53]
  wire  _T_584 = pc_io_read_5_out_bits_way == 2'h2; // @[programmableCache.scala 396:52]
  wire  updateWay_5 = _T_584 & cache_io_cpu_5_resp_valid; // @[programmableCache.scala 396:64]
  wire [2:0] cacheWayWire_5 = {{1'd0}, cache_io_cpu_5_resp_bits_way}; // @[programmableCache.scala 154:28 programmableCache.scala 213:25]
  wire [1:0] pcWire_5_way = pc_io_read_5_out_bits_way; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [2:0] _T_575 = updateWay_5 ? cacheWayWire_5 : {{1'd0}, pcWire_5_way}; // @[programmableCache.scala 386:45]
  wire  firstLineNextRoutine_5 = _GEN_993 == 32'h0; // @[programmableCache.scala 392:72]
  wire [15:0] _T_579 = pcWire_5_pc + 16'h1; // @[programmableCache.scala 393:81]
  wire [15:0] _T_581 = _T_579 + compUnit_5_io_pc; // @[programmableCache.scala 393:87]
  wire [2:0] _T_586 = updateWay_5 ? cacheWayWire_5 : {{1'd0}, pc_io_read_5_out_bits_way}; // @[programmableCache.scala 398:46]
  wire  _T_618 = actionReg_6_io_deq_bits_action_actionType == 4'h0; // @[programmableCache.scala 371:73]
  wire  isCacheAction_6 = _T_618 & actionReg_6_io_deq_valid; // @[programmableCache.scala 371:82]
  wire  _T_620 = actionReg_6_io_deq_bits_action_actionType == 4'h2; // @[programmableCache.scala 372:77]
  wire  _T_624 = actionReg_6_io_deq_bits_action_actionType == 4'h4; // @[programmableCache.scala 374:72]
  wire  _T_626 = actionReg_6_io_deq_bits_action_actionType >= 4'h8; // @[programmableCache.scala 375:73]
  wire [15:0] pcWire_6_pc = pc_io_read_6_out_bits_pc; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [31:0] _GEN_1117 = 6'h1 == pcWire_6_pc[5:0] ? 32'h10000001 : 32'h0; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1118 = 6'h2 == pcWire_6_pc[5:0] ? 32'h34 : _GEN_1117; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1119 = 6'h3 == pcWire_6_pc[5:0] ? 32'hc0000010 : _GEN_1118; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1120 = 6'h4 == pcWire_6_pc[5:0] ? 32'h1000000b : _GEN_1119; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1121 = 6'h5 == pcWire_6_pc[5:0] ? 32'hf0007003 : _GEN_1120; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1122 = 6'h6 == pcWire_6_pc[5:0] ? 32'hf000d013 : _GEN_1121; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1123 = 6'h7 == pcWire_6_pc[5:0] ? 32'h80000405 : _GEN_1122; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1124 = 6'h8 == pcWire_6_pc[5:0] ? 32'hf0015013 : _GEN_1123; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1125 = 6'h9 == pcWire_6_pc[5:0] ? 32'h80000405 : _GEN_1124; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1126 = 6'ha == pcWire_6_pc[5:0] ? 32'h90000005 : _GEN_1125; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1127 = 6'hb == pcWire_6_pc[5:0] ? 32'he07ff011 : _GEN_1126; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1128 = 6'hc == pcWire_6_pc[5:0] ? 32'he06b2016 : _GEN_1127; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1129 = 6'hd == pcWire_6_pc[5:0] ? 32'h10000000 : _GEN_1128; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1130 = 6'he == pcWire_6_pc[5:0] ? 32'he03ff011 : _GEN_1129; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1131 = 6'hf == pcWire_6_pc[5:0] ? 32'he0003404 : _GEN_1130; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1132 = 6'h10 == pcWire_6_pc[5:0] ? 32'hc0000010 : _GEN_1131; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1133 = 6'h11 == pcWire_6_pc[5:0] ? 32'he0800410 : _GEN_1132; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1134 = 6'h12 == pcWire_6_pc[5:0] ? 32'h40000203 : _GEN_1133; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1135 = 6'h13 == pcWire_6_pc[5:0] ? 32'h30000001 : _GEN_1134; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1136 = 6'h14 == pcWire_6_pc[5:0] ? 32'h0 : _GEN_1135; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1137 = 6'h15 == pcWire_6_pc[5:0] ? 32'hc0000037 : _GEN_1136; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1138 = 6'h16 == pcWire_6_pc[5:0] ? 32'h10000000 : _GEN_1137; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1139 = 6'h17 == pcWire_6_pc[5:0] ? 32'h10000002 : _GEN_1138; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1140 = 6'h18 == pcWire_6_pc[5:0] ? 32'h30000000 : _GEN_1139; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1141 = 6'h19 == pcWire_6_pc[5:0] ? 32'h0 : _GEN_1140; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1142 = 6'h1a == pcWire_6_pc[5:0] ? 32'hc0000010 : _GEN_1141; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1143 = 6'h1b == pcWire_6_pc[5:0] ? 32'he0003404 : _GEN_1142; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1144 = 6'h1c == pcWire_6_pc[5:0] ? 32'ha0000010 : _GEN_1143; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1145 = 6'h1d == pcWire_6_pc[5:0] ? 32'h40000203 : _GEN_1144; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1146 = 6'h1e == pcWire_6_pc[5:0] ? 32'h30000002 : _GEN_1145; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1147 = 6'h1f == pcWire_6_pc[5:0] ? 32'h0 : _GEN_1146; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1148 = 6'h20 == pcWire_6_pc[5:0] ? 32'heffff000 : _GEN_1147; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1149 = 6'h21 == pcWire_6_pc[5:0] ? 32'he0010014 : _GEN_1148; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1150 = 6'h22 == pcWire_6_pc[5:0] ? 32'h80001008 : _GEN_1149; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1151 = 6'h23 == pcWire_6_pc[5:0] ? 32'hc0000011 : _GEN_1150; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1152 = 6'h24 == pcWire_6_pc[5:0] ? 32'h90001027 : _GEN_1151; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1153 = 6'h25 == pcWire_6_pc[5:0] ? 32'h10000000 : _GEN_1152; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1154 = 6'h26 == pcWire_6_pc[5:0] ? 32'h80 : _GEN_1153; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1155 = 6'h27 == pcWire_6_pc[5:0] ? 32'h100 : _GEN_1154; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1156 = 6'h28 == pcWire_6_pc[5:0] ? 32'he0020004 : _GEN_1155; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1157 = 6'h29 == pcWire_6_pc[5:0] ? 32'hc0000011 : _GEN_1156; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1158 = 6'h2a == pcWire_6_pc[5:0] ? 32'he0001820 : _GEN_1157; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1159 = 6'h2b == pcWire_6_pc[5:0] ? 32'h80002436 : _GEN_1158; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1160 = 6'h2c == pcWire_6_pc[5:0] ? 32'h10000000 : _GEN_1159; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1161 = 6'h2d == pcWire_6_pc[5:0] ? 32'he001d403 : _GEN_1160; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1162 = 6'h2e == pcWire_6_pc[5:0] ? 32'ha0000010 : _GEN_1161; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1163 = 6'h2f == pcWire_6_pc[5:0] ? 32'h40000203 : _GEN_1162; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1164 = 6'h30 == pcWire_6_pc[5:0] ? 32'h10000002 : _GEN_1163; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1165 = 6'h31 == pcWire_6_pc[5:0] ? 32'h30000003 : _GEN_1164; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1166 = 6'h32 == pcWire_6_pc[5:0] ? 32'h0 : _GEN_1165; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1167 = 6'h33 == pcWire_6_pc[5:0] ? 32'h34 : _GEN_1166; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1168 = 6'h34 == pcWire_6_pc[5:0] ? 32'h80 : _GEN_1167; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1169 = 6'h35 == pcWire_6_pc[5:0] ? 32'h100 : _GEN_1168; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1170 = 6'h36 == pcWire_6_pc[5:0] ? 32'h30000002 : _GEN_1169; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1171 = 6'h37 == pcWire_6_pc[5:0] ? 32'h0 : _GEN_1170; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1172 = 6'h38 == pcWire_6_pc[5:0] ? 32'h30000002 : _GEN_1171; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1173 = 6'h39 == pcWire_6_pc[5:0] ? 32'h0 : _GEN_1172; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1174 = 6'h3a == pcWire_6_pc[5:0] ? 32'h30000003 : _GEN_1173; // @[Gem5CacheLogic.scala 110:53]
  wire  _T_641 = pc_io_read_6_out_bits_way == 2'h2; // @[programmableCache.scala 396:52]
  wire  updateWay_6 = _T_641 & cache_io_cpu_6_resp_valid; // @[programmableCache.scala 396:64]
  wire [2:0] cacheWayWire_6 = {{1'd0}, cache_io_cpu_6_resp_bits_way}; // @[programmableCache.scala 154:28 programmableCache.scala 213:25]
  wire [1:0] pcWire_6_way = pc_io_read_6_out_bits_way; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [2:0] _T_632 = updateWay_6 ? cacheWayWire_6 : {{1'd0}, pcWire_6_way}; // @[programmableCache.scala 386:45]
  wire  firstLineNextRoutine_6 = _GEN_1174 == 32'h0; // @[programmableCache.scala 392:72]
  wire [15:0] _T_636 = pcWire_6_pc + 16'h1; // @[programmableCache.scala 393:81]
  wire [15:0] _T_638 = _T_636 + compUnit_6_io_pc; // @[programmableCache.scala 393:87]
  wire [2:0] _T_643 = updateWay_6 ? cacheWayWire_6 : {{1'd0}, pc_io_read_6_out_bits_way}; // @[programmableCache.scala 398:46]
  wire  _T_675 = actionReg_7_io_deq_bits_action_actionType == 4'h0; // @[programmableCache.scala 371:73]
  wire  isCacheAction_7 = _T_675 & actionReg_7_io_deq_valid; // @[programmableCache.scala 371:82]
  wire  _T_677 = actionReg_7_io_deq_bits_action_actionType == 4'h2; // @[programmableCache.scala 372:77]
  wire  _T_681 = actionReg_7_io_deq_bits_action_actionType == 4'h4; // @[programmableCache.scala 374:72]
  wire  _T_683 = actionReg_7_io_deq_bits_action_actionType >= 4'h8; // @[programmableCache.scala 375:73]
  wire [15:0] pcWire_7_pc = pc_io_read_7_out_bits_pc; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [31:0] _GEN_1298 = 6'h1 == pcWire_7_pc[5:0] ? 32'h10000001 : 32'h0; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1299 = 6'h2 == pcWire_7_pc[5:0] ? 32'h34 : _GEN_1298; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1300 = 6'h3 == pcWire_7_pc[5:0] ? 32'hc0000010 : _GEN_1299; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1301 = 6'h4 == pcWire_7_pc[5:0] ? 32'h1000000b : _GEN_1300; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1302 = 6'h5 == pcWire_7_pc[5:0] ? 32'hf0007003 : _GEN_1301; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1303 = 6'h6 == pcWire_7_pc[5:0] ? 32'hf000d013 : _GEN_1302; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1304 = 6'h7 == pcWire_7_pc[5:0] ? 32'h80000405 : _GEN_1303; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1305 = 6'h8 == pcWire_7_pc[5:0] ? 32'hf0015013 : _GEN_1304; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1306 = 6'h9 == pcWire_7_pc[5:0] ? 32'h80000405 : _GEN_1305; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1307 = 6'ha == pcWire_7_pc[5:0] ? 32'h90000005 : _GEN_1306; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1308 = 6'hb == pcWire_7_pc[5:0] ? 32'he07ff011 : _GEN_1307; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1309 = 6'hc == pcWire_7_pc[5:0] ? 32'he06b2016 : _GEN_1308; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1310 = 6'hd == pcWire_7_pc[5:0] ? 32'h10000000 : _GEN_1309; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1311 = 6'he == pcWire_7_pc[5:0] ? 32'he03ff011 : _GEN_1310; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1312 = 6'hf == pcWire_7_pc[5:0] ? 32'he0003404 : _GEN_1311; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1313 = 6'h10 == pcWire_7_pc[5:0] ? 32'hc0000010 : _GEN_1312; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1314 = 6'h11 == pcWire_7_pc[5:0] ? 32'he0800410 : _GEN_1313; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1315 = 6'h12 == pcWire_7_pc[5:0] ? 32'h40000203 : _GEN_1314; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1316 = 6'h13 == pcWire_7_pc[5:0] ? 32'h30000001 : _GEN_1315; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1317 = 6'h14 == pcWire_7_pc[5:0] ? 32'h0 : _GEN_1316; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1318 = 6'h15 == pcWire_7_pc[5:0] ? 32'hc0000037 : _GEN_1317; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1319 = 6'h16 == pcWire_7_pc[5:0] ? 32'h10000000 : _GEN_1318; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1320 = 6'h17 == pcWire_7_pc[5:0] ? 32'h10000002 : _GEN_1319; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1321 = 6'h18 == pcWire_7_pc[5:0] ? 32'h30000000 : _GEN_1320; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1322 = 6'h19 == pcWire_7_pc[5:0] ? 32'h0 : _GEN_1321; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1323 = 6'h1a == pcWire_7_pc[5:0] ? 32'hc0000010 : _GEN_1322; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1324 = 6'h1b == pcWire_7_pc[5:0] ? 32'he0003404 : _GEN_1323; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1325 = 6'h1c == pcWire_7_pc[5:0] ? 32'ha0000010 : _GEN_1324; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1326 = 6'h1d == pcWire_7_pc[5:0] ? 32'h40000203 : _GEN_1325; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1327 = 6'h1e == pcWire_7_pc[5:0] ? 32'h30000002 : _GEN_1326; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1328 = 6'h1f == pcWire_7_pc[5:0] ? 32'h0 : _GEN_1327; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1329 = 6'h20 == pcWire_7_pc[5:0] ? 32'heffff000 : _GEN_1328; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1330 = 6'h21 == pcWire_7_pc[5:0] ? 32'he0010014 : _GEN_1329; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1331 = 6'h22 == pcWire_7_pc[5:0] ? 32'h80001008 : _GEN_1330; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1332 = 6'h23 == pcWire_7_pc[5:0] ? 32'hc0000011 : _GEN_1331; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1333 = 6'h24 == pcWire_7_pc[5:0] ? 32'h90001027 : _GEN_1332; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1334 = 6'h25 == pcWire_7_pc[5:0] ? 32'h10000000 : _GEN_1333; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1335 = 6'h26 == pcWire_7_pc[5:0] ? 32'h80 : _GEN_1334; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1336 = 6'h27 == pcWire_7_pc[5:0] ? 32'h100 : _GEN_1335; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1337 = 6'h28 == pcWire_7_pc[5:0] ? 32'he0020004 : _GEN_1336; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1338 = 6'h29 == pcWire_7_pc[5:0] ? 32'hc0000011 : _GEN_1337; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1339 = 6'h2a == pcWire_7_pc[5:0] ? 32'he0001820 : _GEN_1338; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1340 = 6'h2b == pcWire_7_pc[5:0] ? 32'h80002436 : _GEN_1339; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1341 = 6'h2c == pcWire_7_pc[5:0] ? 32'h10000000 : _GEN_1340; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1342 = 6'h2d == pcWire_7_pc[5:0] ? 32'he001d403 : _GEN_1341; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1343 = 6'h2e == pcWire_7_pc[5:0] ? 32'ha0000010 : _GEN_1342; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1344 = 6'h2f == pcWire_7_pc[5:0] ? 32'h40000203 : _GEN_1343; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1345 = 6'h30 == pcWire_7_pc[5:0] ? 32'h10000002 : _GEN_1344; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1346 = 6'h31 == pcWire_7_pc[5:0] ? 32'h30000003 : _GEN_1345; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1347 = 6'h32 == pcWire_7_pc[5:0] ? 32'h0 : _GEN_1346; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1348 = 6'h33 == pcWire_7_pc[5:0] ? 32'h34 : _GEN_1347; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1349 = 6'h34 == pcWire_7_pc[5:0] ? 32'h80 : _GEN_1348; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1350 = 6'h35 == pcWire_7_pc[5:0] ? 32'h100 : _GEN_1349; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1351 = 6'h36 == pcWire_7_pc[5:0] ? 32'h30000002 : _GEN_1350; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1352 = 6'h37 == pcWire_7_pc[5:0] ? 32'h0 : _GEN_1351; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1353 = 6'h38 == pcWire_7_pc[5:0] ? 32'h30000002 : _GEN_1352; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1354 = 6'h39 == pcWire_7_pc[5:0] ? 32'h0 : _GEN_1353; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_1355 = 6'h3a == pcWire_7_pc[5:0] ? 32'h30000003 : _GEN_1354; // @[Gem5CacheLogic.scala 110:53]
  wire  _T_698 = pc_io_read_7_out_bits_way == 2'h2; // @[programmableCache.scala 396:52]
  wire  updateWay_7 = _T_698 & cache_io_cpu_7_resp_valid; // @[programmableCache.scala 396:64]
  wire [2:0] cacheWayWire_7 = {{1'd0}, cache_io_cpu_7_resp_bits_way}; // @[programmableCache.scala 154:28 programmableCache.scala 213:25]
  wire [1:0] pcWire_7_way = pc_io_read_7_out_bits_way; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [2:0] _T_689 = updateWay_7 ? cacheWayWire_7 : {{1'd0}, pcWire_7_way}; // @[programmableCache.scala 386:45]
  wire  firstLineNextRoutine_7 = _GEN_1355 == 32'h0; // @[programmableCache.scala 392:72]
  wire [15:0] _T_693 = pcWire_7_pc + 16'h1; // @[programmableCache.scala 393:81]
  wire [15:0] _T_695 = _T_693 + compUnit_7_io_pc; // @[programmableCache.scala 393:87]
  wire [2:0] _T_700 = updateWay_7 ? cacheWayWire_7 : {{1'd0}, pc_io_read_7_out_bits_way}; // @[programmableCache.scala 398:46]
  wire [31:0] instruction_bits_addr = inputArbiter_io_out_bits_addr; // @[programmableCache.scala 110:27 programmableCache.scala 252:17]
  wire  _T_741 = mimoQ_io_deq_bits_0_way != 2'h2; // @[programmableCache.scala 471:83]
  wire [63:0] _GEN_1479 = 2'h1 == actionReg_0_io_deq_bits_action_signals[2:1] ? compUnit_0_io_reg_file_1 : _GEN_207; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1480 = 2'h2 == actionReg_0_io_deq_bits_action_signals[2:1] ? compUnit_0_io_reg_file_2 : _GEN_1479; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1481 = 2'h3 == actionReg_0_io_deq_bits_action_signals[2:1] ? compUnit_0_io_reg_file_3 : _GEN_1480; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1483 = 2'h1 == actionReg_1_io_deq_bits_action_signals[2:1] ? compUnit_1_io_reg_file_1 : _GEN_388; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1484 = 2'h2 == actionReg_1_io_deq_bits_action_signals[2:1] ? compUnit_1_io_reg_file_2 : _GEN_1483; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1485 = 2'h3 == actionReg_1_io_deq_bits_action_signals[2:1] ? compUnit_1_io_reg_file_3 : _GEN_1484; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1487 = 2'h1 == actionReg_2_io_deq_bits_action_signals[2:1] ? compUnit_2_io_reg_file_1 : _GEN_569; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1488 = 2'h2 == actionReg_2_io_deq_bits_action_signals[2:1] ? compUnit_2_io_reg_file_2 : _GEN_1487; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1489 = 2'h3 == actionReg_2_io_deq_bits_action_signals[2:1] ? compUnit_2_io_reg_file_3 : _GEN_1488; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1491 = 2'h1 == actionReg_3_io_deq_bits_action_signals[2:1] ? compUnit_3_io_reg_file_1 : _GEN_750; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1492 = 2'h2 == actionReg_3_io_deq_bits_action_signals[2:1] ? compUnit_3_io_reg_file_2 : _GEN_1491; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1493 = 2'h3 == actionReg_3_io_deq_bits_action_signals[2:1] ? compUnit_3_io_reg_file_3 : _GEN_1492; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1495 = 2'h1 == actionReg_4_io_deq_bits_action_signals[2:1] ? compUnit_4_io_reg_file_1 : _GEN_931; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1496 = 2'h2 == actionReg_4_io_deq_bits_action_signals[2:1] ? compUnit_4_io_reg_file_2 : _GEN_1495; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1497 = 2'h3 == actionReg_4_io_deq_bits_action_signals[2:1] ? compUnit_4_io_reg_file_3 : _GEN_1496; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1499 = 2'h1 == actionReg_5_io_deq_bits_action_signals[2:1] ? compUnit_5_io_reg_file_1 : _GEN_1112; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1500 = 2'h2 == actionReg_5_io_deq_bits_action_signals[2:1] ? compUnit_5_io_reg_file_2 : _GEN_1499; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1501 = 2'h3 == actionReg_5_io_deq_bits_action_signals[2:1] ? compUnit_5_io_reg_file_3 : _GEN_1500; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1503 = 2'h1 == actionReg_6_io_deq_bits_action_signals[2:1] ? compUnit_6_io_reg_file_1 : _GEN_1293; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1504 = 2'h2 == actionReg_6_io_deq_bits_action_signals[2:1] ? compUnit_6_io_reg_file_2 : _GEN_1503; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1505 = 2'h3 == actionReg_6_io_deq_bits_action_signals[2:1] ? compUnit_6_io_reg_file_3 : _GEN_1504; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1507 = 2'h1 == actionReg_7_io_deq_bits_action_signals[2:1] ? compUnit_7_io_reg_file_1 : _GEN_1474; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1508 = 2'h2 == actionReg_7_io_deq_bits_action_signals[2:1] ? compUnit_7_io_reg_file_2 : _GEN_1507; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_1509 = 2'h3 == actionReg_7_io_deq_bits_action_signals[2:1] ? compUnit_7_io_reg_file_3 : _GEN_1508; // @[programmableCache.scala 487:47]
  reg [31:0] _T_783; // @[programmableCache.scala 511:55]
  wire  _T_784 = probeWay_io_deq_ready & probeWay_io_deq_valid; // @[Decoupled.scala 40:37]
  reg [1:0] _T_785; // @[programmableCache.scala 531:49]
  reg [31:0] _T_786; // @[programmableCache.scala 531:90]
  reg [63:0] _T_787; // @[programmableCache.scala 531:138]
  wire  _T_789 = ~reset; // @[programmableCache.scala 531:15]
  reg [1:0] _T_790; // @[programmableCache.scala 532:21]
  wire  _T_791 = _T_790 == 2'h3; // @[programmableCache.scala 532:46]
  reg  _T_798; // @[programmableCache.scala 538:31]
  wire  _T_808 = instruction_ready & instruction_valid; // @[Decoupled.scala 40:37]
  wire  _T_811 = _T_141 & _T_161; // @[programmableCache.scala 557:48]
  wire  _T_814 = _T_141 & _T_158; // @[programmableCache.scala 558:48]
  wire  _T_819 = _T_141 & _T_142; // @[programmableCache.scala 559:48]
  wire  hitLD = _T_153; // @[programmableCache.scala 134:29 programmableCache.scala 276:11]
  wire [2:0] replaceWayInputCache = {{1'd0}, _T_270}; // @[programmableCache.scala 162:36 programmableCache.scala 365:26]
  wire  _GEN_1543 = _T_784 & _T_791; // @[programmableCache.scala 533:19]
  wire  _GEN_1545 = _GEN_1543 & hitLD; // @[programmableCache.scala 535:23]
  wire  _GEN_1547 = ~hitLD; // @[programmableCache.scala 537:23]
  wire  _GEN_1548 = _GEN_1543 & _GEN_1547; // @[programmableCache.scala 537:23]
  wire  _GEN_1549 = _GEN_1548 & isLocked; // @[programmableCache.scala 537:23]
  wire  _GEN_1553 = ~isLocked; // @[programmableCache.scala 539:23]
  wire  _GEN_1554 = _GEN_1548 & _GEN_1553; // @[programmableCache.scala 539:23]
  wire  _GEN_1555 = _GEN_1554 & _T_798; // @[programmableCache.scala 539:23]
  wire  _GEN_1561 = ~_T_798; // @[programmableCache.scala 541:23]
  wire  _GEN_1562 = _GEN_1554 & _GEN_1561; // @[programmableCache.scala 541:23]
  wire  _GEN_1563 = _GEN_1562 & hit; // @[programmableCache.scala 541:23]
  wire  _GEN_1571 = ~hit; // @[programmableCache.scala 543:23]
  wire  _GEN_1572 = _GEN_1562 & _GEN_1571; // @[programmableCache.scala 543:23]
  Gem5Cache cache ( // @[programmableCache.scala 52:26]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_cpu_0_req_valid(cache_io_cpu_0_req_valid),
    .io_cpu_0_req_bits_addr(cache_io_cpu_0_req_bits_addr),
    .io_cpu_0_req_bits_command(cache_io_cpu_0_req_bits_command),
    .io_cpu_0_req_bits_way(cache_io_cpu_0_req_bits_way),
    .io_cpu_0_req_bits_replaceWay(cache_io_cpu_0_req_bits_replaceWay),
    .io_cpu_0_resp_valid(cache_io_cpu_0_resp_valid),
    .io_cpu_0_resp_bits_iswrite(cache_io_cpu_0_resp_bits_iswrite),
    .io_cpu_0_resp_bits_way(cache_io_cpu_0_resp_bits_way),
    .io_cpu_1_req_valid(cache_io_cpu_1_req_valid),
    .io_cpu_1_req_bits_addr(cache_io_cpu_1_req_bits_addr),
    .io_cpu_1_req_bits_command(cache_io_cpu_1_req_bits_command),
    .io_cpu_1_req_bits_way(cache_io_cpu_1_req_bits_way),
    .io_cpu_1_req_bits_replaceWay(cache_io_cpu_1_req_bits_replaceWay),
    .io_cpu_1_resp_valid(cache_io_cpu_1_resp_valid),
    .io_cpu_1_resp_bits_iswrite(cache_io_cpu_1_resp_bits_iswrite),
    .io_cpu_1_resp_bits_way(cache_io_cpu_1_resp_bits_way),
    .io_cpu_2_req_valid(cache_io_cpu_2_req_valid),
    .io_cpu_2_req_bits_addr(cache_io_cpu_2_req_bits_addr),
    .io_cpu_2_req_bits_command(cache_io_cpu_2_req_bits_command),
    .io_cpu_2_req_bits_way(cache_io_cpu_2_req_bits_way),
    .io_cpu_2_req_bits_replaceWay(cache_io_cpu_2_req_bits_replaceWay),
    .io_cpu_2_resp_valid(cache_io_cpu_2_resp_valid),
    .io_cpu_2_resp_bits_iswrite(cache_io_cpu_2_resp_bits_iswrite),
    .io_cpu_2_resp_bits_way(cache_io_cpu_2_resp_bits_way),
    .io_cpu_3_req_valid(cache_io_cpu_3_req_valid),
    .io_cpu_3_req_bits_addr(cache_io_cpu_3_req_bits_addr),
    .io_cpu_3_req_bits_command(cache_io_cpu_3_req_bits_command),
    .io_cpu_3_req_bits_way(cache_io_cpu_3_req_bits_way),
    .io_cpu_3_req_bits_replaceWay(cache_io_cpu_3_req_bits_replaceWay),
    .io_cpu_3_resp_valid(cache_io_cpu_3_resp_valid),
    .io_cpu_3_resp_bits_iswrite(cache_io_cpu_3_resp_bits_iswrite),
    .io_cpu_3_resp_bits_way(cache_io_cpu_3_resp_bits_way),
    .io_cpu_4_req_valid(cache_io_cpu_4_req_valid),
    .io_cpu_4_req_bits_addr(cache_io_cpu_4_req_bits_addr),
    .io_cpu_4_req_bits_command(cache_io_cpu_4_req_bits_command),
    .io_cpu_4_req_bits_way(cache_io_cpu_4_req_bits_way),
    .io_cpu_4_req_bits_replaceWay(cache_io_cpu_4_req_bits_replaceWay),
    .io_cpu_4_resp_valid(cache_io_cpu_4_resp_valid),
    .io_cpu_4_resp_bits_iswrite(cache_io_cpu_4_resp_bits_iswrite),
    .io_cpu_4_resp_bits_way(cache_io_cpu_4_resp_bits_way),
    .io_cpu_5_req_valid(cache_io_cpu_5_req_valid),
    .io_cpu_5_req_bits_addr(cache_io_cpu_5_req_bits_addr),
    .io_cpu_5_req_bits_command(cache_io_cpu_5_req_bits_command),
    .io_cpu_5_req_bits_way(cache_io_cpu_5_req_bits_way),
    .io_cpu_5_req_bits_replaceWay(cache_io_cpu_5_req_bits_replaceWay),
    .io_cpu_5_resp_valid(cache_io_cpu_5_resp_valid),
    .io_cpu_5_resp_bits_iswrite(cache_io_cpu_5_resp_bits_iswrite),
    .io_cpu_5_resp_bits_way(cache_io_cpu_5_resp_bits_way),
    .io_cpu_6_req_valid(cache_io_cpu_6_req_valid),
    .io_cpu_6_req_bits_addr(cache_io_cpu_6_req_bits_addr),
    .io_cpu_6_req_bits_command(cache_io_cpu_6_req_bits_command),
    .io_cpu_6_req_bits_way(cache_io_cpu_6_req_bits_way),
    .io_cpu_6_req_bits_replaceWay(cache_io_cpu_6_req_bits_replaceWay),
    .io_cpu_6_resp_valid(cache_io_cpu_6_resp_valid),
    .io_cpu_6_resp_bits_iswrite(cache_io_cpu_6_resp_bits_iswrite),
    .io_cpu_6_resp_bits_way(cache_io_cpu_6_resp_bits_way),
    .io_cpu_7_req_valid(cache_io_cpu_7_req_valid),
    .io_cpu_7_req_bits_addr(cache_io_cpu_7_req_bits_addr),
    .io_cpu_7_req_bits_data(cache_io_cpu_7_req_bits_data),
    .io_cpu_7_req_bits_command(cache_io_cpu_7_req_bits_command),
    .io_cpu_7_req_bits_way(cache_io_cpu_7_req_bits_way),
    .io_cpu_7_req_bits_replaceWay(cache_io_cpu_7_req_bits_replaceWay),
    .io_cpu_7_resp_valid(cache_io_cpu_7_resp_valid),
    .io_cpu_7_resp_bits_iswrite(cache_io_cpu_7_resp_bits_iswrite),
    .io_cpu_7_resp_bits_way(cache_io_cpu_7_resp_bits_way),
    .io_probe_req_valid(cache_io_probe_req_valid),
    .io_probe_req_bits_addr(cache_io_probe_req_bits_addr),
    .io_probe_req_bits_command(cache_io_probe_req_bits_command),
    .io_probe_resp_valid(cache_io_probe_resp_valid),
    .io_probe_resp_bits_way(cache_io_probe_resp_bits_way),
    .io_probe_multiWay_valid(cache_io_probe_multiWay_valid),
    .io_probe_multiWay_bits_way_0(cache_io_probe_multiWay_bits_way_0),
    .io_probe_multiWay_bits_way_1(cache_io_probe_multiWay_bits_way_1),
    .io_probe_multiWay_bits_addr(cache_io_probe_multiWay_bits_addr),
    .io_bipassLD_in_valid(cache_io_bipassLD_in_valid),
    .io_bipassLD_in_bits_addr(cache_io_bipassLD_in_bits_addr),
    .io_bipassLD_in_bits_way(cache_io_bipassLD_in_bits_way),
    .io_bipassLD_out_valid(cache_io_bipassLD_out_valid),
    .io_bipassLD_out_bits_data(cache_io_bipassLD_out_bits_data)
  );
  TBETable tbe ( // @[programmableCache.scala 53:26]
    .clock(tbe_clock),
    .reset(tbe_reset),
    .io_write_0_valid(tbe_io_write_0_valid),
    .io_write_0_bits_addr(tbe_io_write_0_bits_addr),
    .io_write_0_bits_command(tbe_io_write_0_bits_command),
    .io_write_0_bits_mask(tbe_io_write_0_bits_mask),
    .io_write_0_bits_inputTBE_state_state(tbe_io_write_0_bits_inputTBE_state_state),
    .io_write_0_bits_inputTBE_way(tbe_io_write_0_bits_inputTBE_way),
    .io_write_0_bits_inputTBE_fields_0(tbe_io_write_0_bits_inputTBE_fields_0),
    .io_write_1_valid(tbe_io_write_1_valid),
    .io_write_1_bits_addr(tbe_io_write_1_bits_addr),
    .io_write_1_bits_command(tbe_io_write_1_bits_command),
    .io_write_1_bits_mask(tbe_io_write_1_bits_mask),
    .io_write_1_bits_inputTBE_state_state(tbe_io_write_1_bits_inputTBE_state_state),
    .io_write_1_bits_inputTBE_way(tbe_io_write_1_bits_inputTBE_way),
    .io_write_1_bits_inputTBE_fields_0(tbe_io_write_1_bits_inputTBE_fields_0),
    .io_write_2_valid(tbe_io_write_2_valid),
    .io_write_2_bits_addr(tbe_io_write_2_bits_addr),
    .io_write_2_bits_command(tbe_io_write_2_bits_command),
    .io_write_2_bits_mask(tbe_io_write_2_bits_mask),
    .io_write_2_bits_inputTBE_state_state(tbe_io_write_2_bits_inputTBE_state_state),
    .io_write_2_bits_inputTBE_way(tbe_io_write_2_bits_inputTBE_way),
    .io_write_2_bits_inputTBE_fields_0(tbe_io_write_2_bits_inputTBE_fields_0),
    .io_write_3_valid(tbe_io_write_3_valid),
    .io_write_3_bits_addr(tbe_io_write_3_bits_addr),
    .io_write_3_bits_command(tbe_io_write_3_bits_command),
    .io_write_3_bits_mask(tbe_io_write_3_bits_mask),
    .io_write_3_bits_inputTBE_state_state(tbe_io_write_3_bits_inputTBE_state_state),
    .io_write_3_bits_inputTBE_way(tbe_io_write_3_bits_inputTBE_way),
    .io_write_3_bits_inputTBE_fields_0(tbe_io_write_3_bits_inputTBE_fields_0),
    .io_write_4_valid(tbe_io_write_4_valid),
    .io_write_4_bits_addr(tbe_io_write_4_bits_addr),
    .io_write_4_bits_command(tbe_io_write_4_bits_command),
    .io_write_4_bits_mask(tbe_io_write_4_bits_mask),
    .io_write_4_bits_inputTBE_state_state(tbe_io_write_4_bits_inputTBE_state_state),
    .io_write_4_bits_inputTBE_way(tbe_io_write_4_bits_inputTBE_way),
    .io_write_4_bits_inputTBE_fields_0(tbe_io_write_4_bits_inputTBE_fields_0),
    .io_write_5_valid(tbe_io_write_5_valid),
    .io_write_5_bits_addr(tbe_io_write_5_bits_addr),
    .io_write_5_bits_command(tbe_io_write_5_bits_command),
    .io_write_5_bits_mask(tbe_io_write_5_bits_mask),
    .io_write_5_bits_inputTBE_state_state(tbe_io_write_5_bits_inputTBE_state_state),
    .io_write_5_bits_inputTBE_way(tbe_io_write_5_bits_inputTBE_way),
    .io_write_5_bits_inputTBE_fields_0(tbe_io_write_5_bits_inputTBE_fields_0),
    .io_write_6_valid(tbe_io_write_6_valid),
    .io_write_6_bits_addr(tbe_io_write_6_bits_addr),
    .io_write_6_bits_command(tbe_io_write_6_bits_command),
    .io_write_6_bits_mask(tbe_io_write_6_bits_mask),
    .io_write_6_bits_inputTBE_state_state(tbe_io_write_6_bits_inputTBE_state_state),
    .io_write_6_bits_inputTBE_way(tbe_io_write_6_bits_inputTBE_way),
    .io_write_6_bits_inputTBE_fields_0(tbe_io_write_6_bits_inputTBE_fields_0),
    .io_write_7_valid(tbe_io_write_7_valid),
    .io_write_7_bits_addr(tbe_io_write_7_bits_addr),
    .io_write_7_bits_command(tbe_io_write_7_bits_command),
    .io_write_7_bits_mask(tbe_io_write_7_bits_mask),
    .io_write_7_bits_inputTBE_state_state(tbe_io_write_7_bits_inputTBE_state_state),
    .io_write_7_bits_inputTBE_way(tbe_io_write_7_bits_inputTBE_way),
    .io_write_7_bits_inputTBE_fields_0(tbe_io_write_7_bits_inputTBE_fields_0),
    .io_read_valid(tbe_io_read_valid),
    .io_read_bits_addr(tbe_io_read_bits_addr),
    .io_outputTBE_bits_state_state(tbe_io_outputTBE_bits_state_state),
    .io_outputTBE_bits_way(tbe_io_outputTBE_bits_way),
    .io_outputTBE_bits_fields_0(tbe_io_outputTBE_bits_fields_0),
    .io_isFull(tbe_io_isFull)
  );
  lockVector lockMem ( // @[programmableCache.scala 54:26]
    .clock(lockMem_clock),
    .reset(lockMem_reset),
    .io_lock_in_valid(lockMem_io_lock_in_valid),
    .io_lock_in_bits_addr(lockMem_io_lock_in_bits_addr),
    .io_probe_out_valid(lockMem_io_probe_out_valid),
    .io_probe_out_bits(lockMem_io_probe_out_bits),
    .io_probe_in_valid(lockMem_io_probe_in_valid),
    .io_probe_in_bits_addr(lockMem_io_probe_in_bits_addr),
    .io_unLock_0_in_valid(lockMem_io_unLock_0_in_valid),
    .io_unLock_0_in_bits_addr(lockMem_io_unLock_0_in_bits_addr),
    .io_unLock_1_in_valid(lockMem_io_unLock_1_in_valid),
    .io_unLock_1_in_bits_addr(lockMem_io_unLock_1_in_bits_addr),
    .io_unLock_2_in_valid(lockMem_io_unLock_2_in_valid),
    .io_unLock_2_in_bits_addr(lockMem_io_unLock_2_in_bits_addr),
    .io_unLock_3_in_valid(lockMem_io_unLock_3_in_valid),
    .io_unLock_3_in_bits_addr(lockMem_io_unLock_3_in_bits_addr),
    .io_unLock_4_in_valid(lockMem_io_unLock_4_in_valid),
    .io_unLock_4_in_bits_addr(lockMem_io_unLock_4_in_bits_addr),
    .io_unLock_5_in_valid(lockMem_io_unLock_5_in_valid),
    .io_unLock_5_in_bits_addr(lockMem_io_unLock_5_in_bits_addr),
    .io_unLock_6_in_valid(lockMem_io_unLock_6_in_valid),
    .io_unLock_6_in_bits_addr(lockMem_io_unLock_6_in_bits_addr),
    .io_unLock_7_in_valid(lockMem_io_unLock_7_in_valid),
    .io_unLock_7_in_bits_addr(lockMem_io_unLock_7_in_bits_addr)
  );
  stateMem stateMem ( // @[programmableCache.scala 55:27]
    .clock(stateMem_clock),
    .reset(stateMem_reset),
    .io_in_0_valid(stateMem_io_in_0_valid),
    .io_in_0_bits_state_state(stateMem_io_in_0_bits_state_state),
    .io_in_0_bits_addr(stateMem_io_in_0_bits_addr),
    .io_in_0_bits_way(stateMem_io_in_0_bits_way),
    .io_in_1_valid(stateMem_io_in_1_valid),
    .io_in_1_bits_state_state(stateMem_io_in_1_bits_state_state),
    .io_in_1_bits_addr(stateMem_io_in_1_bits_addr),
    .io_in_1_bits_way(stateMem_io_in_1_bits_way),
    .io_in_2_valid(stateMem_io_in_2_valid),
    .io_in_2_bits_state_state(stateMem_io_in_2_bits_state_state),
    .io_in_2_bits_addr(stateMem_io_in_2_bits_addr),
    .io_in_2_bits_way(stateMem_io_in_2_bits_way),
    .io_in_3_valid(stateMem_io_in_3_valid),
    .io_in_3_bits_state_state(stateMem_io_in_3_bits_state_state),
    .io_in_3_bits_addr(stateMem_io_in_3_bits_addr),
    .io_in_3_bits_way(stateMem_io_in_3_bits_way),
    .io_in_4_valid(stateMem_io_in_4_valid),
    .io_in_4_bits_state_state(stateMem_io_in_4_bits_state_state),
    .io_in_4_bits_addr(stateMem_io_in_4_bits_addr),
    .io_in_4_bits_way(stateMem_io_in_4_bits_way),
    .io_in_5_valid(stateMem_io_in_5_valid),
    .io_in_5_bits_state_state(stateMem_io_in_5_bits_state_state),
    .io_in_5_bits_addr(stateMem_io_in_5_bits_addr),
    .io_in_5_bits_way(stateMem_io_in_5_bits_way),
    .io_in_6_valid(stateMem_io_in_6_valid),
    .io_in_6_bits_state_state(stateMem_io_in_6_bits_state_state),
    .io_in_6_bits_addr(stateMem_io_in_6_bits_addr),
    .io_in_6_bits_way(stateMem_io_in_6_bits_way),
    .io_in_7_valid(stateMem_io_in_7_valid),
    .io_in_7_bits_state_state(stateMem_io_in_7_bits_state_state),
    .io_in_7_bits_addr(stateMem_io_in_7_bits_addr),
    .io_in_7_bits_way(stateMem_io_in_7_bits_way),
    .io_in_8_valid(stateMem_io_in_8_valid),
    .io_in_8_bits_addr(stateMem_io_in_8_bits_addr),
    .io_in_8_bits_way(stateMem_io_in_8_bits_way),
    .io_out_valid(stateMem_io_out_valid),
    .io_out_bits_state(stateMem_io_out_bits_state)
  );
  PC pc ( // @[programmableCache.scala 56:26]
    .clock(pc_clock),
    .reset(pc_reset),
    .io_write_ready(pc_io_write_ready),
    .io_write_valid(pc_io_write_valid),
    .io_write_bits_addr(pc_io_write_bits_addr),
    .io_write_bits_way(pc_io_write_bits_way),
    .io_write_bits_data(pc_io_write_bits_data),
    .io_write_bits_replaceWay(pc_io_write_bits_replaceWay),
    .io_write_bits_tbeFields_0(pc_io_write_bits_tbeFields_0),
    .io_write_bits_pc(pc_io_write_bits_pc),
    .io_read_0_in_bits_data_way(pc_io_read_0_in_bits_data_way),
    .io_read_0_in_bits_data_pc(pc_io_read_0_in_bits_data_pc),
    .io_read_0_in_bits_data_valid(pc_io_read_0_in_bits_data_valid),
    .io_read_0_out_bits_addr(pc_io_read_0_out_bits_addr),
    .io_read_0_out_bits_way(pc_io_read_0_out_bits_way),
    .io_read_0_out_bits_data(pc_io_read_0_out_bits_data),
    .io_read_0_out_bits_replaceWay(pc_io_read_0_out_bits_replaceWay),
    .io_read_0_out_bits_tbeFields_0(pc_io_read_0_out_bits_tbeFields_0),
    .io_read_0_out_bits_pc(pc_io_read_0_out_bits_pc),
    .io_read_0_out_bits_valid(pc_io_read_0_out_bits_valid),
    .io_read_1_in_bits_data_way(pc_io_read_1_in_bits_data_way),
    .io_read_1_in_bits_data_pc(pc_io_read_1_in_bits_data_pc),
    .io_read_1_in_bits_data_valid(pc_io_read_1_in_bits_data_valid),
    .io_read_1_out_bits_addr(pc_io_read_1_out_bits_addr),
    .io_read_1_out_bits_way(pc_io_read_1_out_bits_way),
    .io_read_1_out_bits_data(pc_io_read_1_out_bits_data),
    .io_read_1_out_bits_replaceWay(pc_io_read_1_out_bits_replaceWay),
    .io_read_1_out_bits_tbeFields_0(pc_io_read_1_out_bits_tbeFields_0),
    .io_read_1_out_bits_pc(pc_io_read_1_out_bits_pc),
    .io_read_1_out_bits_valid(pc_io_read_1_out_bits_valid),
    .io_read_2_in_bits_data_way(pc_io_read_2_in_bits_data_way),
    .io_read_2_in_bits_data_pc(pc_io_read_2_in_bits_data_pc),
    .io_read_2_in_bits_data_valid(pc_io_read_2_in_bits_data_valid),
    .io_read_2_out_bits_addr(pc_io_read_2_out_bits_addr),
    .io_read_2_out_bits_way(pc_io_read_2_out_bits_way),
    .io_read_2_out_bits_data(pc_io_read_2_out_bits_data),
    .io_read_2_out_bits_replaceWay(pc_io_read_2_out_bits_replaceWay),
    .io_read_2_out_bits_tbeFields_0(pc_io_read_2_out_bits_tbeFields_0),
    .io_read_2_out_bits_pc(pc_io_read_2_out_bits_pc),
    .io_read_2_out_bits_valid(pc_io_read_2_out_bits_valid),
    .io_read_3_in_bits_data_way(pc_io_read_3_in_bits_data_way),
    .io_read_3_in_bits_data_pc(pc_io_read_3_in_bits_data_pc),
    .io_read_3_in_bits_data_valid(pc_io_read_3_in_bits_data_valid),
    .io_read_3_out_bits_addr(pc_io_read_3_out_bits_addr),
    .io_read_3_out_bits_way(pc_io_read_3_out_bits_way),
    .io_read_3_out_bits_data(pc_io_read_3_out_bits_data),
    .io_read_3_out_bits_replaceWay(pc_io_read_3_out_bits_replaceWay),
    .io_read_3_out_bits_tbeFields_0(pc_io_read_3_out_bits_tbeFields_0),
    .io_read_3_out_bits_pc(pc_io_read_3_out_bits_pc),
    .io_read_3_out_bits_valid(pc_io_read_3_out_bits_valid),
    .io_read_4_in_bits_data_way(pc_io_read_4_in_bits_data_way),
    .io_read_4_in_bits_data_pc(pc_io_read_4_in_bits_data_pc),
    .io_read_4_in_bits_data_valid(pc_io_read_4_in_bits_data_valid),
    .io_read_4_out_bits_addr(pc_io_read_4_out_bits_addr),
    .io_read_4_out_bits_way(pc_io_read_4_out_bits_way),
    .io_read_4_out_bits_data(pc_io_read_4_out_bits_data),
    .io_read_4_out_bits_replaceWay(pc_io_read_4_out_bits_replaceWay),
    .io_read_4_out_bits_tbeFields_0(pc_io_read_4_out_bits_tbeFields_0),
    .io_read_4_out_bits_pc(pc_io_read_4_out_bits_pc),
    .io_read_4_out_bits_valid(pc_io_read_4_out_bits_valid),
    .io_read_5_in_bits_data_way(pc_io_read_5_in_bits_data_way),
    .io_read_5_in_bits_data_pc(pc_io_read_5_in_bits_data_pc),
    .io_read_5_in_bits_data_valid(pc_io_read_5_in_bits_data_valid),
    .io_read_5_out_bits_addr(pc_io_read_5_out_bits_addr),
    .io_read_5_out_bits_way(pc_io_read_5_out_bits_way),
    .io_read_5_out_bits_data(pc_io_read_5_out_bits_data),
    .io_read_5_out_bits_replaceWay(pc_io_read_5_out_bits_replaceWay),
    .io_read_5_out_bits_tbeFields_0(pc_io_read_5_out_bits_tbeFields_0),
    .io_read_5_out_bits_pc(pc_io_read_5_out_bits_pc),
    .io_read_5_out_bits_valid(pc_io_read_5_out_bits_valid),
    .io_read_6_in_bits_data_way(pc_io_read_6_in_bits_data_way),
    .io_read_6_in_bits_data_pc(pc_io_read_6_in_bits_data_pc),
    .io_read_6_in_bits_data_valid(pc_io_read_6_in_bits_data_valid),
    .io_read_6_out_bits_addr(pc_io_read_6_out_bits_addr),
    .io_read_6_out_bits_way(pc_io_read_6_out_bits_way),
    .io_read_6_out_bits_data(pc_io_read_6_out_bits_data),
    .io_read_6_out_bits_replaceWay(pc_io_read_6_out_bits_replaceWay),
    .io_read_6_out_bits_tbeFields_0(pc_io_read_6_out_bits_tbeFields_0),
    .io_read_6_out_bits_pc(pc_io_read_6_out_bits_pc),
    .io_read_6_out_bits_valid(pc_io_read_6_out_bits_valid),
    .io_read_7_in_bits_data_way(pc_io_read_7_in_bits_data_way),
    .io_read_7_in_bits_data_pc(pc_io_read_7_in_bits_data_pc),
    .io_read_7_in_bits_data_valid(pc_io_read_7_in_bits_data_valid),
    .io_read_7_out_bits_addr(pc_io_read_7_out_bits_addr),
    .io_read_7_out_bits_way(pc_io_read_7_out_bits_way),
    .io_read_7_out_bits_data(pc_io_read_7_out_bits_data),
    .io_read_7_out_bits_replaceWay(pc_io_read_7_out_bits_replaceWay),
    .io_read_7_out_bits_tbeFields_0(pc_io_read_7_out_bits_tbeFields_0),
    .io_read_7_out_bits_pc(pc_io_read_7_out_bits_pc),
    .io_read_7_out_bits_valid(pc_io_read_7_out_bits_valid),
    .io_isFull(pc_io_isFull)
  );
  Arbiter_3 inputArbiter ( // @[programmableCache.scala 57:33]
    .io_in_0_valid(inputArbiter_io_in_0_valid),
    .io_in_0_bits_event(inputArbiter_io_in_0_bits_event),
    .io_in_0_bits_addr(inputArbiter_io_in_0_bits_addr),
    .io_in_0_bits_data(inputArbiter_io_in_0_bits_data),
    .io_in_1_ready(inputArbiter_io_in_1_ready),
    .io_in_1_valid(inputArbiter_io_in_1_valid),
    .io_in_1_bits_event(inputArbiter_io_in_1_bits_event),
    .io_in_1_bits_addr(inputArbiter_io_in_1_bits_addr),
    .io_in_1_bits_data(inputArbiter_io_in_1_bits_data),
    .io_in_2_valid(inputArbiter_io_in_2_valid),
    .io_in_2_bits_event(inputArbiter_io_in_2_bits_event),
    .io_in_2_bits_addr(inputArbiter_io_in_2_bits_addr),
    .io_in_2_bits_data(inputArbiter_io_in_2_bits_data),
    .io_in_3_valid(inputArbiter_io_in_3_valid),
    .io_in_3_bits_event(inputArbiter_io_in_3_bits_event),
    .io_in_3_bits_addr(inputArbiter_io_in_3_bits_addr),
    .io_in_3_bits_data(inputArbiter_io_in_3_bits_data),
    .io_out_ready(inputArbiter_io_out_ready),
    .io_out_valid(inputArbiter_io_out_valid),
    .io_out_bits_event(inputArbiter_io_out_bits_event),
    .io_out_bits_addr(inputArbiter_io_out_bits_addr),
    .io_out_bits_data(inputArbiter_io_out_bits_data),
    .io_chosen(inputArbiter_io_chosen)
  );
  RRArbiter_2 outReqArbiter ( // @[programmableCache.scala 58:33]
    .clock(outReqArbiter_clock),
    .io_in_0_ready(outReqArbiter_io_in_0_ready),
    .io_in_0_valid(outReqArbiter_io_in_0_valid),
    .io_in_0_bits_req_addr(outReqArbiter_io_in_0_bits_req_addr),
    .io_in_0_bits_req_inst(outReqArbiter_io_in_0_bits_req_inst),
    .io_in_0_bits_req_data(outReqArbiter_io_in_0_bits_req_data),
    .io_in_1_ready(outReqArbiter_io_in_1_ready),
    .io_in_1_valid(outReqArbiter_io_in_1_valid),
    .io_in_1_bits_req_addr(outReqArbiter_io_in_1_bits_req_addr),
    .io_in_1_bits_req_inst(outReqArbiter_io_in_1_bits_req_inst),
    .io_in_1_bits_req_data(outReqArbiter_io_in_1_bits_req_data),
    .io_in_2_ready(outReqArbiter_io_in_2_ready),
    .io_in_2_valid(outReqArbiter_io_in_2_valid),
    .io_in_2_bits_req_addr(outReqArbiter_io_in_2_bits_req_addr),
    .io_in_2_bits_req_inst(outReqArbiter_io_in_2_bits_req_inst),
    .io_in_2_bits_req_data(outReqArbiter_io_in_2_bits_req_data),
    .io_in_3_ready(outReqArbiter_io_in_3_ready),
    .io_in_3_valid(outReqArbiter_io_in_3_valid),
    .io_in_3_bits_req_addr(outReqArbiter_io_in_3_bits_req_addr),
    .io_in_3_bits_req_inst(outReqArbiter_io_in_3_bits_req_inst),
    .io_in_3_bits_req_data(outReqArbiter_io_in_3_bits_req_data),
    .io_in_4_ready(outReqArbiter_io_in_4_ready),
    .io_in_4_valid(outReqArbiter_io_in_4_valid),
    .io_in_4_bits_req_addr(outReqArbiter_io_in_4_bits_req_addr),
    .io_in_4_bits_req_inst(outReqArbiter_io_in_4_bits_req_inst),
    .io_in_4_bits_req_data(outReqArbiter_io_in_4_bits_req_data),
    .io_in_5_ready(outReqArbiter_io_in_5_ready),
    .io_in_5_valid(outReqArbiter_io_in_5_valid),
    .io_in_5_bits_req_addr(outReqArbiter_io_in_5_bits_req_addr),
    .io_in_5_bits_req_inst(outReqArbiter_io_in_5_bits_req_inst),
    .io_in_5_bits_req_data(outReqArbiter_io_in_5_bits_req_data),
    .io_in_6_ready(outReqArbiter_io_in_6_ready),
    .io_in_6_valid(outReqArbiter_io_in_6_valid),
    .io_in_6_bits_req_addr(outReqArbiter_io_in_6_bits_req_addr),
    .io_in_6_bits_req_inst(outReqArbiter_io_in_6_bits_req_inst),
    .io_in_6_bits_req_data(outReqArbiter_io_in_6_bits_req_data),
    .io_in_7_ready(outReqArbiter_io_in_7_ready),
    .io_in_7_valid(outReqArbiter_io_in_7_valid),
    .io_in_7_bits_req_addr(outReqArbiter_io_in_7_bits_req_addr),
    .io_in_7_bits_req_inst(outReqArbiter_io_in_7_bits_req_inst),
    .io_in_7_bits_req_data(outReqArbiter_io_in_7_bits_req_data),
    .io_out_valid(outReqArbiter_io_out_valid),
    .io_out_bits_req_addr(outReqArbiter_io_out_bits_req_addr),
    .io_out_bits_req_inst(outReqArbiter_io_out_bits_req_inst),
    .io_out_bits_req_data(outReqArbiter_io_out_bits_req_data),
    .io_chosen(outReqArbiter_io_chosen)
  );
  Arbiter_4 outRespArbiter ( // @[programmableCache.scala 59:33]
    .io_in_0_valid(outRespArbiter_io_in_0_valid),
    .io_in_0_bits_addr(outRespArbiter_io_in_0_bits_addr),
    .io_in_1_valid(outRespArbiter_io_in_1_valid),
    .io_in_1_bits_addr(outRespArbiter_io_in_1_bits_addr),
    .io_in_2_valid(outRespArbiter_io_in_2_valid),
    .io_in_2_bits_addr(outRespArbiter_io_in_2_bits_addr),
    .io_in_3_valid(outRespArbiter_io_in_3_valid),
    .io_in_3_bits_addr(outRespArbiter_io_in_3_bits_addr),
    .io_in_4_valid(outRespArbiter_io_in_4_valid),
    .io_in_4_bits_addr(outRespArbiter_io_in_4_bits_addr),
    .io_in_5_valid(outRespArbiter_io_in_5_valid),
    .io_in_5_bits_addr(outRespArbiter_io_in_5_bits_addr),
    .io_in_6_valid(outRespArbiter_io_in_6_valid),
    .io_in_6_bits_addr(outRespArbiter_io_in_6_bits_addr),
    .io_in_7_valid(outRespArbiter_io_in_7_valid),
    .io_in_7_bits_addr(outRespArbiter_io_in_7_bits_addr),
    .io_in_8_valid(outRespArbiter_io_in_8_valid),
    .io_in_8_bits_addr(outRespArbiter_io_in_8_bits_addr),
    .io_out_valid(outRespArbiter_io_out_valid),
    .io_out_bits_addr(outRespArbiter_io_out_bits_addr)
  );
  Arbiter_5 feedbackArbiter ( // @[programmableCache.scala 60:34]
    .io_in_0_ready(feedbackArbiter_io_in_0_ready),
    .io_in_0_valid(feedbackArbiter_io_in_0_valid),
    .io_in_0_bits_event(feedbackArbiter_io_in_0_bits_event),
    .io_in_0_bits_addr(feedbackArbiter_io_in_0_bits_addr),
    .io_in_0_bits_data(feedbackArbiter_io_in_0_bits_data),
    .io_in_1_ready(feedbackArbiter_io_in_1_ready),
    .io_in_1_valid(feedbackArbiter_io_in_1_valid),
    .io_in_1_bits_event(feedbackArbiter_io_in_1_bits_event),
    .io_in_1_bits_addr(feedbackArbiter_io_in_1_bits_addr),
    .io_in_1_bits_data(feedbackArbiter_io_in_1_bits_data),
    .io_in_2_ready(feedbackArbiter_io_in_2_ready),
    .io_in_2_valid(feedbackArbiter_io_in_2_valid),
    .io_in_2_bits_event(feedbackArbiter_io_in_2_bits_event),
    .io_in_2_bits_addr(feedbackArbiter_io_in_2_bits_addr),
    .io_in_2_bits_data(feedbackArbiter_io_in_2_bits_data),
    .io_in_3_ready(feedbackArbiter_io_in_3_ready),
    .io_in_3_valid(feedbackArbiter_io_in_3_valid),
    .io_in_3_bits_event(feedbackArbiter_io_in_3_bits_event),
    .io_in_3_bits_addr(feedbackArbiter_io_in_3_bits_addr),
    .io_in_3_bits_data(feedbackArbiter_io_in_3_bits_data),
    .io_in_4_ready(feedbackArbiter_io_in_4_ready),
    .io_in_4_valid(feedbackArbiter_io_in_4_valid),
    .io_in_4_bits_event(feedbackArbiter_io_in_4_bits_event),
    .io_in_4_bits_addr(feedbackArbiter_io_in_4_bits_addr),
    .io_in_4_bits_data(feedbackArbiter_io_in_4_bits_data),
    .io_in_5_ready(feedbackArbiter_io_in_5_ready),
    .io_in_5_valid(feedbackArbiter_io_in_5_valid),
    .io_in_5_bits_event(feedbackArbiter_io_in_5_bits_event),
    .io_in_5_bits_addr(feedbackArbiter_io_in_5_bits_addr),
    .io_in_5_bits_data(feedbackArbiter_io_in_5_bits_data),
    .io_in_6_ready(feedbackArbiter_io_in_6_ready),
    .io_in_6_valid(feedbackArbiter_io_in_6_valid),
    .io_in_6_bits_event(feedbackArbiter_io_in_6_bits_event),
    .io_in_6_bits_addr(feedbackArbiter_io_in_6_bits_addr),
    .io_in_6_bits_data(feedbackArbiter_io_in_6_bits_data),
    .io_in_7_ready(feedbackArbiter_io_in_7_ready),
    .io_in_7_valid(feedbackArbiter_io_in_7_valid),
    .io_in_7_bits_event(feedbackArbiter_io_in_7_bits_event),
    .io_in_7_bits_addr(feedbackArbiter_io_in_7_bits_addr),
    .io_in_7_bits_data(feedbackArbiter_io_in_7_bits_data),
    .io_out_ready(feedbackArbiter_io_out_ready),
    .io_out_valid(feedbackArbiter_io_out_valid),
    .io_out_bits_event(feedbackArbiter_io_out_bits_event),
    .io_out_bits_addr(feedbackArbiter_io_out_bits_addr),
    .io_out_bits_data(feedbackArbiter_io_out_bits_data)
  );
  Queue_7 input_ ( // @[programmableCache.scala 90:23]
    .clock(input__clock),
    .reset(input__reset),
    .io_enq_ready(input__io_enq_ready),
    .io_enq_valid(input__io_enq_valid),
    .io_enq_bits_inst_event(input__io_enq_bits_inst_event),
    .io_enq_bits_inst_addr(input__io_enq_bits_inst_addr),
    .io_enq_bits_inst_data(input__io_enq_bits_inst_data),
    .io_enq_bits_tbeOut_state_state(input__io_enq_bits_tbeOut_state_state),
    .io_enq_bits_tbeOut_way(input__io_enq_bits_tbeOut_way),
    .io_enq_bits_tbeOut_fields_0(input__io_enq_bits_tbeOut_fields_0),
    .io_deq_ready(input__io_deq_ready),
    .io_deq_valid(input__io_deq_valid),
    .io_deq_bits_inst_event(input__io_deq_bits_inst_event),
    .io_deq_bits_inst_addr(input__io_deq_bits_inst_addr),
    .io_deq_bits_inst_data(input__io_deq_bits_inst_data),
    .io_deq_bits_tbeOut_state_state(input__io_deq_bits_tbeOut_state_state),
    .io_deq_bits_tbeOut_way(input__io_deq_bits_tbeOut_way),
    .io_deq_bits_tbeOut_fields_0(input__io_deq_bits_tbeOut_fields_0)
  );
  Queue_8 respPortQueue_0 ( // @[programmableCache.scala 93:27]
    .clock(respPortQueue_0_clock),
    .reset(respPortQueue_0_reset),
    .io_enq_ready(respPortQueue_0_io_enq_ready),
    .io_enq_valid(respPortQueue_0_io_enq_valid),
    .io_enq_bits_event(respPortQueue_0_io_enq_bits_event),
    .io_enq_bits_addr(respPortQueue_0_io_enq_bits_addr),
    .io_enq_bits_data(respPortQueue_0_io_enq_bits_data),
    .io_deq_ready(respPortQueue_0_io_deq_ready),
    .io_deq_valid(respPortQueue_0_io_deq_valid),
    .io_deq_bits_event(respPortQueue_0_io_deq_bits_event),
    .io_deq_bits_addr(respPortQueue_0_io_deq_bits_addr),
    .io_deq_bits_data(respPortQueue_0_io_deq_bits_data)
  );
  Queue_8 respPortQueue_1 ( // @[programmableCache.scala 93:27]
    .clock(respPortQueue_1_clock),
    .reset(respPortQueue_1_reset),
    .io_enq_ready(respPortQueue_1_io_enq_ready),
    .io_enq_valid(respPortQueue_1_io_enq_valid),
    .io_enq_bits_event(respPortQueue_1_io_enq_bits_event),
    .io_enq_bits_addr(respPortQueue_1_io_enq_bits_addr),
    .io_enq_bits_data(respPortQueue_1_io_enq_bits_data),
    .io_deq_ready(respPortQueue_1_io_deq_ready),
    .io_deq_valid(respPortQueue_1_io_deq_valid),
    .io_deq_bits_event(respPortQueue_1_io_deq_bits_event),
    .io_deq_bits_addr(respPortQueue_1_io_deq_bits_addr),
    .io_deq_bits_data(respPortQueue_1_io_deq_bits_data)
  );
  Queue_8 respPortQueue_2 ( // @[programmableCache.scala 93:27]
    .clock(respPortQueue_2_clock),
    .reset(respPortQueue_2_reset),
    .io_enq_ready(respPortQueue_2_io_enq_ready),
    .io_enq_valid(respPortQueue_2_io_enq_valid),
    .io_enq_bits_event(respPortQueue_2_io_enq_bits_event),
    .io_enq_bits_addr(respPortQueue_2_io_enq_bits_addr),
    .io_enq_bits_data(respPortQueue_2_io_enq_bits_data),
    .io_deq_ready(respPortQueue_2_io_deq_ready),
    .io_deq_valid(respPortQueue_2_io_deq_valid),
    .io_deq_bits_event(respPortQueue_2_io_deq_bits_event),
    .io_deq_bits_addr(respPortQueue_2_io_deq_bits_addr),
    .io_deq_bits_data(respPortQueue_2_io_deq_bits_data)
  );
  Queue_8 respPortQueue_3 ( // @[programmableCache.scala 93:27]
    .clock(respPortQueue_3_clock),
    .reset(respPortQueue_3_reset),
    .io_enq_ready(respPortQueue_3_io_enq_ready),
    .io_enq_valid(respPortQueue_3_io_enq_valid),
    .io_enq_bits_event(respPortQueue_3_io_enq_bits_event),
    .io_enq_bits_addr(respPortQueue_3_io_enq_bits_addr),
    .io_enq_bits_data(respPortQueue_3_io_enq_bits_data),
    .io_deq_ready(respPortQueue_3_io_deq_ready),
    .io_deq_valid(respPortQueue_3_io_deq_valid),
    .io_deq_bits_event(respPortQueue_3_io_deq_bits_event),
    .io_deq_bits_addr(respPortQueue_3_io_deq_bits_addr),
    .io_deq_bits_data(respPortQueue_3_io_deq_bits_data)
  );
  Queue_8 respPortQueue_4 ( // @[programmableCache.scala 93:27]
    .clock(respPortQueue_4_clock),
    .reset(respPortQueue_4_reset),
    .io_enq_ready(respPortQueue_4_io_enq_ready),
    .io_enq_valid(respPortQueue_4_io_enq_valid),
    .io_enq_bits_event(respPortQueue_4_io_enq_bits_event),
    .io_enq_bits_addr(respPortQueue_4_io_enq_bits_addr),
    .io_enq_bits_data(respPortQueue_4_io_enq_bits_data),
    .io_deq_ready(respPortQueue_4_io_deq_ready),
    .io_deq_valid(respPortQueue_4_io_deq_valid),
    .io_deq_bits_event(respPortQueue_4_io_deq_bits_event),
    .io_deq_bits_addr(respPortQueue_4_io_deq_bits_addr),
    .io_deq_bits_data(respPortQueue_4_io_deq_bits_data)
  );
  Queue_8 respPortQueue_5 ( // @[programmableCache.scala 93:27]
    .clock(respPortQueue_5_clock),
    .reset(respPortQueue_5_reset),
    .io_enq_ready(respPortQueue_5_io_enq_ready),
    .io_enq_valid(respPortQueue_5_io_enq_valid),
    .io_enq_bits_event(respPortQueue_5_io_enq_bits_event),
    .io_enq_bits_addr(respPortQueue_5_io_enq_bits_addr),
    .io_enq_bits_data(respPortQueue_5_io_enq_bits_data),
    .io_deq_ready(respPortQueue_5_io_deq_ready),
    .io_deq_valid(respPortQueue_5_io_deq_valid),
    .io_deq_bits_event(respPortQueue_5_io_deq_bits_event),
    .io_deq_bits_addr(respPortQueue_5_io_deq_bits_addr),
    .io_deq_bits_data(respPortQueue_5_io_deq_bits_data)
  );
  Queue_8 respPortQueue_6 ( // @[programmableCache.scala 93:27]
    .clock(respPortQueue_6_clock),
    .reset(respPortQueue_6_reset),
    .io_enq_ready(respPortQueue_6_io_enq_ready),
    .io_enq_valid(respPortQueue_6_io_enq_valid),
    .io_enq_bits_event(respPortQueue_6_io_enq_bits_event),
    .io_enq_bits_addr(respPortQueue_6_io_enq_bits_addr),
    .io_enq_bits_data(respPortQueue_6_io_enq_bits_data),
    .io_deq_ready(respPortQueue_6_io_deq_ready),
    .io_deq_valid(respPortQueue_6_io_deq_valid),
    .io_deq_bits_event(respPortQueue_6_io_deq_bits_event),
    .io_deq_bits_addr(respPortQueue_6_io_deq_bits_addr),
    .io_deq_bits_data(respPortQueue_6_io_deq_bits_data)
  );
  Queue_8 respPortQueue_7 ( // @[programmableCache.scala 93:27]
    .clock(respPortQueue_7_clock),
    .reset(respPortQueue_7_reset),
    .io_enq_ready(respPortQueue_7_io_enq_ready),
    .io_enq_valid(respPortQueue_7_io_enq_valid),
    .io_enq_bits_event(respPortQueue_7_io_enq_bits_event),
    .io_enq_bits_addr(respPortQueue_7_io_enq_bits_addr),
    .io_enq_bits_data(respPortQueue_7_io_enq_bits_data),
    .io_deq_ready(respPortQueue_7_io_deq_ready),
    .io_deq_valid(respPortQueue_7_io_deq_valid),
    .io_deq_bits_event(respPortQueue_7_io_deq_bits_event),
    .io_deq_bits_addr(respPortQueue_7_io_deq_bits_addr),
    .io_deq_bits_data(respPortQueue_7_io_deq_bits_data)
  );
  Queue_8 respPortQueue_8 ( // @[programmableCache.scala 93:27]
    .clock(respPortQueue_8_clock),
    .reset(respPortQueue_8_reset),
    .io_enq_ready(respPortQueue_8_io_enq_ready),
    .io_enq_valid(respPortQueue_8_io_enq_valid),
    .io_enq_bits_event(respPortQueue_8_io_enq_bits_event),
    .io_enq_bits_addr(respPortQueue_8_io_enq_bits_addr),
    .io_enq_bits_data(respPortQueue_8_io_enq_bits_data),
    .io_deq_ready(respPortQueue_8_io_deq_ready),
    .io_deq_valid(respPortQueue_8_io_deq_valid),
    .io_deq_bits_event(respPortQueue_8_io_deq_bits_event),
    .io_deq_bits_addr(respPortQueue_8_io_deq_bits_addr),
    .io_deq_bits_data(respPortQueue_8_io_deq_bits_data)
  );
  Queue_17 reqPortQueue_0 ( // @[programmableCache.scala 98:27]
    .clock(reqPortQueue_0_clock),
    .reset(reqPortQueue_0_reset),
    .io_enq_ready(reqPortQueue_0_io_enq_ready),
    .io_enq_valid(reqPortQueue_0_io_enq_valid),
    .io_enq_bits_addr(reqPortQueue_0_io_enq_bits_addr),
    .io_enq_bits_inst(reqPortQueue_0_io_enq_bits_inst),
    .io_enq_bits_data(reqPortQueue_0_io_enq_bits_data),
    .io_deq_ready(reqPortQueue_0_io_deq_ready),
    .io_deq_valid(reqPortQueue_0_io_deq_valid),
    .io_deq_bits_addr(reqPortQueue_0_io_deq_bits_addr),
    .io_deq_bits_inst(reqPortQueue_0_io_deq_bits_inst),
    .io_deq_bits_data(reqPortQueue_0_io_deq_bits_data)
  );
  Queue_17 reqPortQueue_1 ( // @[programmableCache.scala 98:27]
    .clock(reqPortQueue_1_clock),
    .reset(reqPortQueue_1_reset),
    .io_enq_ready(reqPortQueue_1_io_enq_ready),
    .io_enq_valid(reqPortQueue_1_io_enq_valid),
    .io_enq_bits_addr(reqPortQueue_1_io_enq_bits_addr),
    .io_enq_bits_inst(reqPortQueue_1_io_enq_bits_inst),
    .io_enq_bits_data(reqPortQueue_1_io_enq_bits_data),
    .io_deq_ready(reqPortQueue_1_io_deq_ready),
    .io_deq_valid(reqPortQueue_1_io_deq_valid),
    .io_deq_bits_addr(reqPortQueue_1_io_deq_bits_addr),
    .io_deq_bits_inst(reqPortQueue_1_io_deq_bits_inst),
    .io_deq_bits_data(reqPortQueue_1_io_deq_bits_data)
  );
  Queue_17 reqPortQueue_2 ( // @[programmableCache.scala 98:27]
    .clock(reqPortQueue_2_clock),
    .reset(reqPortQueue_2_reset),
    .io_enq_ready(reqPortQueue_2_io_enq_ready),
    .io_enq_valid(reqPortQueue_2_io_enq_valid),
    .io_enq_bits_addr(reqPortQueue_2_io_enq_bits_addr),
    .io_enq_bits_inst(reqPortQueue_2_io_enq_bits_inst),
    .io_enq_bits_data(reqPortQueue_2_io_enq_bits_data),
    .io_deq_ready(reqPortQueue_2_io_deq_ready),
    .io_deq_valid(reqPortQueue_2_io_deq_valid),
    .io_deq_bits_addr(reqPortQueue_2_io_deq_bits_addr),
    .io_deq_bits_inst(reqPortQueue_2_io_deq_bits_inst),
    .io_deq_bits_data(reqPortQueue_2_io_deq_bits_data)
  );
  Queue_17 reqPortQueue_3 ( // @[programmableCache.scala 98:27]
    .clock(reqPortQueue_3_clock),
    .reset(reqPortQueue_3_reset),
    .io_enq_ready(reqPortQueue_3_io_enq_ready),
    .io_enq_valid(reqPortQueue_3_io_enq_valid),
    .io_enq_bits_addr(reqPortQueue_3_io_enq_bits_addr),
    .io_enq_bits_inst(reqPortQueue_3_io_enq_bits_inst),
    .io_enq_bits_data(reqPortQueue_3_io_enq_bits_data),
    .io_deq_ready(reqPortQueue_3_io_deq_ready),
    .io_deq_valid(reqPortQueue_3_io_deq_valid),
    .io_deq_bits_addr(reqPortQueue_3_io_deq_bits_addr),
    .io_deq_bits_inst(reqPortQueue_3_io_deq_bits_inst),
    .io_deq_bits_data(reqPortQueue_3_io_deq_bits_data)
  );
  Queue_17 reqPortQueue_4 ( // @[programmableCache.scala 98:27]
    .clock(reqPortQueue_4_clock),
    .reset(reqPortQueue_4_reset),
    .io_enq_ready(reqPortQueue_4_io_enq_ready),
    .io_enq_valid(reqPortQueue_4_io_enq_valid),
    .io_enq_bits_addr(reqPortQueue_4_io_enq_bits_addr),
    .io_enq_bits_inst(reqPortQueue_4_io_enq_bits_inst),
    .io_enq_bits_data(reqPortQueue_4_io_enq_bits_data),
    .io_deq_ready(reqPortQueue_4_io_deq_ready),
    .io_deq_valid(reqPortQueue_4_io_deq_valid),
    .io_deq_bits_addr(reqPortQueue_4_io_deq_bits_addr),
    .io_deq_bits_inst(reqPortQueue_4_io_deq_bits_inst),
    .io_deq_bits_data(reqPortQueue_4_io_deq_bits_data)
  );
  Queue_17 reqPortQueue_5 ( // @[programmableCache.scala 98:27]
    .clock(reqPortQueue_5_clock),
    .reset(reqPortQueue_5_reset),
    .io_enq_ready(reqPortQueue_5_io_enq_ready),
    .io_enq_valid(reqPortQueue_5_io_enq_valid),
    .io_enq_bits_addr(reqPortQueue_5_io_enq_bits_addr),
    .io_enq_bits_inst(reqPortQueue_5_io_enq_bits_inst),
    .io_enq_bits_data(reqPortQueue_5_io_enq_bits_data),
    .io_deq_ready(reqPortQueue_5_io_deq_ready),
    .io_deq_valid(reqPortQueue_5_io_deq_valid),
    .io_deq_bits_addr(reqPortQueue_5_io_deq_bits_addr),
    .io_deq_bits_inst(reqPortQueue_5_io_deq_bits_inst),
    .io_deq_bits_data(reqPortQueue_5_io_deq_bits_data)
  );
  Queue_17 reqPortQueue_6 ( // @[programmableCache.scala 98:27]
    .clock(reqPortQueue_6_clock),
    .reset(reqPortQueue_6_reset),
    .io_enq_ready(reqPortQueue_6_io_enq_ready),
    .io_enq_valid(reqPortQueue_6_io_enq_valid),
    .io_enq_bits_addr(reqPortQueue_6_io_enq_bits_addr),
    .io_enq_bits_inst(reqPortQueue_6_io_enq_bits_inst),
    .io_enq_bits_data(reqPortQueue_6_io_enq_bits_data),
    .io_deq_ready(reqPortQueue_6_io_deq_ready),
    .io_deq_valid(reqPortQueue_6_io_deq_valid),
    .io_deq_bits_addr(reqPortQueue_6_io_deq_bits_addr),
    .io_deq_bits_inst(reqPortQueue_6_io_deq_bits_inst),
    .io_deq_bits_data(reqPortQueue_6_io_deq_bits_data)
  );
  Queue_17 reqPortQueue_7 ( // @[programmableCache.scala 98:27]
    .clock(reqPortQueue_7_clock),
    .reset(reqPortQueue_7_reset),
    .io_enq_ready(reqPortQueue_7_io_enq_ready),
    .io_enq_valid(reqPortQueue_7_io_enq_valid),
    .io_enq_bits_addr(reqPortQueue_7_io_enq_bits_addr),
    .io_enq_bits_inst(reqPortQueue_7_io_enq_bits_inst),
    .io_enq_bits_data(reqPortQueue_7_io_enq_bits_data),
    .io_deq_ready(reqPortQueue_7_io_deq_ready),
    .io_deq_valid(reqPortQueue_7_io_deq_valid),
    .io_deq_bits_addr(reqPortQueue_7_io_deq_bits_addr),
    .io_deq_bits_inst(reqPortQueue_7_io_deq_bits_inst),
    .io_deq_bits_data(reqPortQueue_7_io_deq_bits_data)
  );
  Queue_8 feedbackInQueue_0 ( // @[programmableCache.scala 104:27]
    .clock(feedbackInQueue_0_clock),
    .reset(feedbackInQueue_0_reset),
    .io_enq_ready(feedbackInQueue_0_io_enq_ready),
    .io_enq_valid(feedbackInQueue_0_io_enq_valid),
    .io_enq_bits_event(feedbackInQueue_0_io_enq_bits_event),
    .io_enq_bits_addr(feedbackInQueue_0_io_enq_bits_addr),
    .io_enq_bits_data(feedbackInQueue_0_io_enq_bits_data),
    .io_deq_ready(feedbackInQueue_0_io_deq_ready),
    .io_deq_valid(feedbackInQueue_0_io_deq_valid),
    .io_deq_bits_event(feedbackInQueue_0_io_deq_bits_event),
    .io_deq_bits_addr(feedbackInQueue_0_io_deq_bits_addr),
    .io_deq_bits_data(feedbackInQueue_0_io_deq_bits_data)
  );
  Queue_8 feedbackInQueue_1 ( // @[programmableCache.scala 104:27]
    .clock(feedbackInQueue_1_clock),
    .reset(feedbackInQueue_1_reset),
    .io_enq_ready(feedbackInQueue_1_io_enq_ready),
    .io_enq_valid(feedbackInQueue_1_io_enq_valid),
    .io_enq_bits_event(feedbackInQueue_1_io_enq_bits_event),
    .io_enq_bits_addr(feedbackInQueue_1_io_enq_bits_addr),
    .io_enq_bits_data(feedbackInQueue_1_io_enq_bits_data),
    .io_deq_ready(feedbackInQueue_1_io_deq_ready),
    .io_deq_valid(feedbackInQueue_1_io_deq_valid),
    .io_deq_bits_event(feedbackInQueue_1_io_deq_bits_event),
    .io_deq_bits_addr(feedbackInQueue_1_io_deq_bits_addr),
    .io_deq_bits_data(feedbackInQueue_1_io_deq_bits_data)
  );
  Queue_8 feedbackInQueue_2 ( // @[programmableCache.scala 104:27]
    .clock(feedbackInQueue_2_clock),
    .reset(feedbackInQueue_2_reset),
    .io_enq_ready(feedbackInQueue_2_io_enq_ready),
    .io_enq_valid(feedbackInQueue_2_io_enq_valid),
    .io_enq_bits_event(feedbackInQueue_2_io_enq_bits_event),
    .io_enq_bits_addr(feedbackInQueue_2_io_enq_bits_addr),
    .io_enq_bits_data(feedbackInQueue_2_io_enq_bits_data),
    .io_deq_ready(feedbackInQueue_2_io_deq_ready),
    .io_deq_valid(feedbackInQueue_2_io_deq_valid),
    .io_deq_bits_event(feedbackInQueue_2_io_deq_bits_event),
    .io_deq_bits_addr(feedbackInQueue_2_io_deq_bits_addr),
    .io_deq_bits_data(feedbackInQueue_2_io_deq_bits_data)
  );
  Queue_8 feedbackInQueue_3 ( // @[programmableCache.scala 104:27]
    .clock(feedbackInQueue_3_clock),
    .reset(feedbackInQueue_3_reset),
    .io_enq_ready(feedbackInQueue_3_io_enq_ready),
    .io_enq_valid(feedbackInQueue_3_io_enq_valid),
    .io_enq_bits_event(feedbackInQueue_3_io_enq_bits_event),
    .io_enq_bits_addr(feedbackInQueue_3_io_enq_bits_addr),
    .io_enq_bits_data(feedbackInQueue_3_io_enq_bits_data),
    .io_deq_ready(feedbackInQueue_3_io_deq_ready),
    .io_deq_valid(feedbackInQueue_3_io_deq_valid),
    .io_deq_bits_event(feedbackInQueue_3_io_deq_bits_event),
    .io_deq_bits_addr(feedbackInQueue_3_io_deq_bits_addr),
    .io_deq_bits_data(feedbackInQueue_3_io_deq_bits_data)
  );
  Queue_8 feedbackInQueue_4 ( // @[programmableCache.scala 104:27]
    .clock(feedbackInQueue_4_clock),
    .reset(feedbackInQueue_4_reset),
    .io_enq_ready(feedbackInQueue_4_io_enq_ready),
    .io_enq_valid(feedbackInQueue_4_io_enq_valid),
    .io_enq_bits_event(feedbackInQueue_4_io_enq_bits_event),
    .io_enq_bits_addr(feedbackInQueue_4_io_enq_bits_addr),
    .io_enq_bits_data(feedbackInQueue_4_io_enq_bits_data),
    .io_deq_ready(feedbackInQueue_4_io_deq_ready),
    .io_deq_valid(feedbackInQueue_4_io_deq_valid),
    .io_deq_bits_event(feedbackInQueue_4_io_deq_bits_event),
    .io_deq_bits_addr(feedbackInQueue_4_io_deq_bits_addr),
    .io_deq_bits_data(feedbackInQueue_4_io_deq_bits_data)
  );
  Queue_8 feedbackInQueue_5 ( // @[programmableCache.scala 104:27]
    .clock(feedbackInQueue_5_clock),
    .reset(feedbackInQueue_5_reset),
    .io_enq_ready(feedbackInQueue_5_io_enq_ready),
    .io_enq_valid(feedbackInQueue_5_io_enq_valid),
    .io_enq_bits_event(feedbackInQueue_5_io_enq_bits_event),
    .io_enq_bits_addr(feedbackInQueue_5_io_enq_bits_addr),
    .io_enq_bits_data(feedbackInQueue_5_io_enq_bits_data),
    .io_deq_ready(feedbackInQueue_5_io_deq_ready),
    .io_deq_valid(feedbackInQueue_5_io_deq_valid),
    .io_deq_bits_event(feedbackInQueue_5_io_deq_bits_event),
    .io_deq_bits_addr(feedbackInQueue_5_io_deq_bits_addr),
    .io_deq_bits_data(feedbackInQueue_5_io_deq_bits_data)
  );
  Queue_8 feedbackInQueue_6 ( // @[programmableCache.scala 104:27]
    .clock(feedbackInQueue_6_clock),
    .reset(feedbackInQueue_6_reset),
    .io_enq_ready(feedbackInQueue_6_io_enq_ready),
    .io_enq_valid(feedbackInQueue_6_io_enq_valid),
    .io_enq_bits_event(feedbackInQueue_6_io_enq_bits_event),
    .io_enq_bits_addr(feedbackInQueue_6_io_enq_bits_addr),
    .io_enq_bits_data(feedbackInQueue_6_io_enq_bits_data),
    .io_deq_ready(feedbackInQueue_6_io_deq_ready),
    .io_deq_valid(feedbackInQueue_6_io_deq_valid),
    .io_deq_bits_event(feedbackInQueue_6_io_deq_bits_event),
    .io_deq_bits_addr(feedbackInQueue_6_io_deq_bits_addr),
    .io_deq_bits_data(feedbackInQueue_6_io_deq_bits_data)
  );
  Queue_8 feedbackInQueue_7 ( // @[programmableCache.scala 104:27]
    .clock(feedbackInQueue_7_clock),
    .reset(feedbackInQueue_7_reset),
    .io_enq_ready(feedbackInQueue_7_io_enq_ready),
    .io_enq_valid(feedbackInQueue_7_io_enq_valid),
    .io_enq_bits_event(feedbackInQueue_7_io_enq_bits_event),
    .io_enq_bits_addr(feedbackInQueue_7_io_enq_bits_addr),
    .io_enq_bits_data(feedbackInQueue_7_io_enq_bits_data),
    .io_deq_ready(feedbackInQueue_7_io_deq_ready),
    .io_deq_valid(feedbackInQueue_7_io_deq_valid),
    .io_deq_bits_event(feedbackInQueue_7_io_deq_bits_event),
    .io_deq_bits_addr(feedbackInQueue_7_io_deq_bits_addr),
    .io_deq_bits_data(feedbackInQueue_7_io_deq_bits_data)
  );
  Queue_33 probeWay ( // @[programmableCache.scala 108:26]
    .clock(probeWay_clock),
    .reset(probeWay_reset),
    .io_enq_ready(probeWay_io_enq_ready),
    .io_enq_valid(probeWay_io_enq_valid),
    .io_enq_bits(probeWay_io_enq_bits),
    .io_deq_ready(probeWay_io_deq_ready),
    .io_deq_valid(probeWay_io_deq_valid),
    .io_deq_bits(probeWay_io_deq_bits)
  );
  Queue_8 feedbackOutQueue ( // @[programmableCache.scala 165:34]
    .clock(feedbackOutQueue_clock),
    .reset(feedbackOutQueue_reset),
    .io_enq_ready(feedbackOutQueue_io_enq_ready),
    .io_enq_valid(feedbackOutQueue_io_enq_valid),
    .io_enq_bits_event(feedbackOutQueue_io_enq_bits_event),
    .io_enq_bits_addr(feedbackOutQueue_io_enq_bits_addr),
    .io_enq_bits_data(feedbackOutQueue_io_enq_bits_data),
    .io_deq_ready(feedbackOutQueue_io_deq_ready),
    .io_deq_valid(feedbackOutQueue_io_deq_valid),
    .io_deq_bits_event(feedbackOutQueue_io_deq_bits_event),
    .io_deq_bits_addr(feedbackOutQueue_io_deq_bits_addr),
    .io_deq_bits_data(feedbackOutQueue_io_deq_bits_data)
  );
  Queue_35 routineQueue ( // @[programmableCache.scala 166:30]
    .clock(routineQueue_clock),
    .reset(routineQueue_reset),
    .io_enq_ready(routineQueue_io_enq_ready),
    .io_enq_valid(routineQueue_io_enq_valid),
    .io_enq_bits(routineQueue_io_enq_bits),
    .io_deq_ready(routineQueue_io_deq_ready),
    .io_deq_valid(routineQueue_io_deq_valid),
    .io_deq_bits(routineQueue_io_deq_bits)
  );
  Queue_36 actionReg_0 ( // @[programmableCache.scala 169:32]
    .clock(actionReg_0_clock),
    .reset(actionReg_0_reset),
    .io_enq_ready(actionReg_0_io_enq_ready),
    .io_enq_valid(actionReg_0_io_enq_valid),
    .io_enq_bits_addr(actionReg_0_io_enq_bits_addr),
    .io_enq_bits_way(actionReg_0_io_enq_bits_way),
    .io_enq_bits_data(actionReg_0_io_enq_bits_data),
    .io_enq_bits_replaceWay(actionReg_0_io_enq_bits_replaceWay),
    .io_enq_bits_tbeFields_0(actionReg_0_io_enq_bits_tbeFields_0),
    .io_enq_bits_action_signals(actionReg_0_io_enq_bits_action_signals),
    .io_enq_bits_action_actionType(actionReg_0_io_enq_bits_action_actionType),
    .io_deq_ready(actionReg_0_io_deq_ready),
    .io_deq_valid(actionReg_0_io_deq_valid),
    .io_deq_bits_addr(actionReg_0_io_deq_bits_addr),
    .io_deq_bits_way(actionReg_0_io_deq_bits_way),
    .io_deq_bits_data(actionReg_0_io_deq_bits_data),
    .io_deq_bits_replaceWay(actionReg_0_io_deq_bits_replaceWay),
    .io_deq_bits_tbeFields_0(actionReg_0_io_deq_bits_tbeFields_0),
    .io_deq_bits_action_signals(actionReg_0_io_deq_bits_action_signals),
    .io_deq_bits_action_actionType(actionReg_0_io_deq_bits_action_actionType)
  );
  Queue_36 actionReg_1 ( // @[programmableCache.scala 169:32]
    .clock(actionReg_1_clock),
    .reset(actionReg_1_reset),
    .io_enq_ready(actionReg_1_io_enq_ready),
    .io_enq_valid(actionReg_1_io_enq_valid),
    .io_enq_bits_addr(actionReg_1_io_enq_bits_addr),
    .io_enq_bits_way(actionReg_1_io_enq_bits_way),
    .io_enq_bits_data(actionReg_1_io_enq_bits_data),
    .io_enq_bits_replaceWay(actionReg_1_io_enq_bits_replaceWay),
    .io_enq_bits_tbeFields_0(actionReg_1_io_enq_bits_tbeFields_0),
    .io_enq_bits_action_signals(actionReg_1_io_enq_bits_action_signals),
    .io_enq_bits_action_actionType(actionReg_1_io_enq_bits_action_actionType),
    .io_deq_ready(actionReg_1_io_deq_ready),
    .io_deq_valid(actionReg_1_io_deq_valid),
    .io_deq_bits_addr(actionReg_1_io_deq_bits_addr),
    .io_deq_bits_way(actionReg_1_io_deq_bits_way),
    .io_deq_bits_data(actionReg_1_io_deq_bits_data),
    .io_deq_bits_replaceWay(actionReg_1_io_deq_bits_replaceWay),
    .io_deq_bits_tbeFields_0(actionReg_1_io_deq_bits_tbeFields_0),
    .io_deq_bits_action_signals(actionReg_1_io_deq_bits_action_signals),
    .io_deq_bits_action_actionType(actionReg_1_io_deq_bits_action_actionType)
  );
  Queue_36 actionReg_2 ( // @[programmableCache.scala 169:32]
    .clock(actionReg_2_clock),
    .reset(actionReg_2_reset),
    .io_enq_ready(actionReg_2_io_enq_ready),
    .io_enq_valid(actionReg_2_io_enq_valid),
    .io_enq_bits_addr(actionReg_2_io_enq_bits_addr),
    .io_enq_bits_way(actionReg_2_io_enq_bits_way),
    .io_enq_bits_data(actionReg_2_io_enq_bits_data),
    .io_enq_bits_replaceWay(actionReg_2_io_enq_bits_replaceWay),
    .io_enq_bits_tbeFields_0(actionReg_2_io_enq_bits_tbeFields_0),
    .io_enq_bits_action_signals(actionReg_2_io_enq_bits_action_signals),
    .io_enq_bits_action_actionType(actionReg_2_io_enq_bits_action_actionType),
    .io_deq_ready(actionReg_2_io_deq_ready),
    .io_deq_valid(actionReg_2_io_deq_valid),
    .io_deq_bits_addr(actionReg_2_io_deq_bits_addr),
    .io_deq_bits_way(actionReg_2_io_deq_bits_way),
    .io_deq_bits_data(actionReg_2_io_deq_bits_data),
    .io_deq_bits_replaceWay(actionReg_2_io_deq_bits_replaceWay),
    .io_deq_bits_tbeFields_0(actionReg_2_io_deq_bits_tbeFields_0),
    .io_deq_bits_action_signals(actionReg_2_io_deq_bits_action_signals),
    .io_deq_bits_action_actionType(actionReg_2_io_deq_bits_action_actionType)
  );
  Queue_36 actionReg_3 ( // @[programmableCache.scala 169:32]
    .clock(actionReg_3_clock),
    .reset(actionReg_3_reset),
    .io_enq_ready(actionReg_3_io_enq_ready),
    .io_enq_valid(actionReg_3_io_enq_valid),
    .io_enq_bits_addr(actionReg_3_io_enq_bits_addr),
    .io_enq_bits_way(actionReg_3_io_enq_bits_way),
    .io_enq_bits_data(actionReg_3_io_enq_bits_data),
    .io_enq_bits_replaceWay(actionReg_3_io_enq_bits_replaceWay),
    .io_enq_bits_tbeFields_0(actionReg_3_io_enq_bits_tbeFields_0),
    .io_enq_bits_action_signals(actionReg_3_io_enq_bits_action_signals),
    .io_enq_bits_action_actionType(actionReg_3_io_enq_bits_action_actionType),
    .io_deq_ready(actionReg_3_io_deq_ready),
    .io_deq_valid(actionReg_3_io_deq_valid),
    .io_deq_bits_addr(actionReg_3_io_deq_bits_addr),
    .io_deq_bits_way(actionReg_3_io_deq_bits_way),
    .io_deq_bits_data(actionReg_3_io_deq_bits_data),
    .io_deq_bits_replaceWay(actionReg_3_io_deq_bits_replaceWay),
    .io_deq_bits_tbeFields_0(actionReg_3_io_deq_bits_tbeFields_0),
    .io_deq_bits_action_signals(actionReg_3_io_deq_bits_action_signals),
    .io_deq_bits_action_actionType(actionReg_3_io_deq_bits_action_actionType)
  );
  Queue_36 actionReg_4 ( // @[programmableCache.scala 169:32]
    .clock(actionReg_4_clock),
    .reset(actionReg_4_reset),
    .io_enq_ready(actionReg_4_io_enq_ready),
    .io_enq_valid(actionReg_4_io_enq_valid),
    .io_enq_bits_addr(actionReg_4_io_enq_bits_addr),
    .io_enq_bits_way(actionReg_4_io_enq_bits_way),
    .io_enq_bits_data(actionReg_4_io_enq_bits_data),
    .io_enq_bits_replaceWay(actionReg_4_io_enq_bits_replaceWay),
    .io_enq_bits_tbeFields_0(actionReg_4_io_enq_bits_tbeFields_0),
    .io_enq_bits_action_signals(actionReg_4_io_enq_bits_action_signals),
    .io_enq_bits_action_actionType(actionReg_4_io_enq_bits_action_actionType),
    .io_deq_ready(actionReg_4_io_deq_ready),
    .io_deq_valid(actionReg_4_io_deq_valid),
    .io_deq_bits_addr(actionReg_4_io_deq_bits_addr),
    .io_deq_bits_way(actionReg_4_io_deq_bits_way),
    .io_deq_bits_data(actionReg_4_io_deq_bits_data),
    .io_deq_bits_replaceWay(actionReg_4_io_deq_bits_replaceWay),
    .io_deq_bits_tbeFields_0(actionReg_4_io_deq_bits_tbeFields_0),
    .io_deq_bits_action_signals(actionReg_4_io_deq_bits_action_signals),
    .io_deq_bits_action_actionType(actionReg_4_io_deq_bits_action_actionType)
  );
  Queue_36 actionReg_5 ( // @[programmableCache.scala 169:32]
    .clock(actionReg_5_clock),
    .reset(actionReg_5_reset),
    .io_enq_ready(actionReg_5_io_enq_ready),
    .io_enq_valid(actionReg_5_io_enq_valid),
    .io_enq_bits_addr(actionReg_5_io_enq_bits_addr),
    .io_enq_bits_way(actionReg_5_io_enq_bits_way),
    .io_enq_bits_data(actionReg_5_io_enq_bits_data),
    .io_enq_bits_replaceWay(actionReg_5_io_enq_bits_replaceWay),
    .io_enq_bits_tbeFields_0(actionReg_5_io_enq_bits_tbeFields_0),
    .io_enq_bits_action_signals(actionReg_5_io_enq_bits_action_signals),
    .io_enq_bits_action_actionType(actionReg_5_io_enq_bits_action_actionType),
    .io_deq_ready(actionReg_5_io_deq_ready),
    .io_deq_valid(actionReg_5_io_deq_valid),
    .io_deq_bits_addr(actionReg_5_io_deq_bits_addr),
    .io_deq_bits_way(actionReg_5_io_deq_bits_way),
    .io_deq_bits_data(actionReg_5_io_deq_bits_data),
    .io_deq_bits_replaceWay(actionReg_5_io_deq_bits_replaceWay),
    .io_deq_bits_tbeFields_0(actionReg_5_io_deq_bits_tbeFields_0),
    .io_deq_bits_action_signals(actionReg_5_io_deq_bits_action_signals),
    .io_deq_bits_action_actionType(actionReg_5_io_deq_bits_action_actionType)
  );
  Queue_36 actionReg_6 ( // @[programmableCache.scala 169:32]
    .clock(actionReg_6_clock),
    .reset(actionReg_6_reset),
    .io_enq_ready(actionReg_6_io_enq_ready),
    .io_enq_valid(actionReg_6_io_enq_valid),
    .io_enq_bits_addr(actionReg_6_io_enq_bits_addr),
    .io_enq_bits_way(actionReg_6_io_enq_bits_way),
    .io_enq_bits_data(actionReg_6_io_enq_bits_data),
    .io_enq_bits_replaceWay(actionReg_6_io_enq_bits_replaceWay),
    .io_enq_bits_tbeFields_0(actionReg_6_io_enq_bits_tbeFields_0),
    .io_enq_bits_action_signals(actionReg_6_io_enq_bits_action_signals),
    .io_enq_bits_action_actionType(actionReg_6_io_enq_bits_action_actionType),
    .io_deq_ready(actionReg_6_io_deq_ready),
    .io_deq_valid(actionReg_6_io_deq_valid),
    .io_deq_bits_addr(actionReg_6_io_deq_bits_addr),
    .io_deq_bits_way(actionReg_6_io_deq_bits_way),
    .io_deq_bits_data(actionReg_6_io_deq_bits_data),
    .io_deq_bits_replaceWay(actionReg_6_io_deq_bits_replaceWay),
    .io_deq_bits_tbeFields_0(actionReg_6_io_deq_bits_tbeFields_0),
    .io_deq_bits_action_signals(actionReg_6_io_deq_bits_action_signals),
    .io_deq_bits_action_actionType(actionReg_6_io_deq_bits_action_actionType)
  );
  Queue_36 actionReg_7 ( // @[programmableCache.scala 169:32]
    .clock(actionReg_7_clock),
    .reset(actionReg_7_reset),
    .io_enq_ready(actionReg_7_io_enq_ready),
    .io_enq_valid(actionReg_7_io_enq_valid),
    .io_enq_bits_addr(actionReg_7_io_enq_bits_addr),
    .io_enq_bits_way(actionReg_7_io_enq_bits_way),
    .io_enq_bits_data(actionReg_7_io_enq_bits_data),
    .io_enq_bits_replaceWay(actionReg_7_io_enq_bits_replaceWay),
    .io_enq_bits_tbeFields_0(actionReg_7_io_enq_bits_tbeFields_0),
    .io_enq_bits_action_signals(actionReg_7_io_enq_bits_action_signals),
    .io_enq_bits_action_actionType(actionReg_7_io_enq_bits_action_actionType),
    .io_deq_ready(actionReg_7_io_deq_ready),
    .io_deq_valid(actionReg_7_io_deq_valid),
    .io_deq_bits_addr(actionReg_7_io_deq_bits_addr),
    .io_deq_bits_way(actionReg_7_io_deq_bits_way),
    .io_deq_bits_data(actionReg_7_io_deq_bits_data),
    .io_deq_bits_replaceWay(actionReg_7_io_deq_bits_replaceWay),
    .io_deq_bits_tbeFields_0(actionReg_7_io_deq_bits_tbeFields_0),
    .io_deq_bits_action_signals(actionReg_7_io_deq_bits_action_signals),
    .io_deq_bits_action_actionType(actionReg_7_io_deq_bits_action_actionType)
  );
  MIMOQueue mimoQ ( // @[programmableCache.scala 173:24]
    .clock(mimoQ_clock),
    .reset(mimoQ_reset),
    .io_enq_ready(mimoQ_io_enq_ready),
    .io_enq_valid(mimoQ_io_enq_valid),
    .io_enq_bits_0_way(mimoQ_io_enq_bits_0_way),
    .io_enq_bits_0_addr(mimoQ_io_enq_bits_0_addr),
    .io_enq_bits_1_way(mimoQ_io_enq_bits_1_way),
    .io_enq_bits_1_addr(mimoQ_io_enq_bits_1_addr),
    .io_deq_valid(mimoQ_io_deq_valid),
    .io_deq_bits_0_way(mimoQ_io_deq_bits_0_way),
    .io_deq_bits_0_addr(mimoQ_io_deq_bits_0_addr),
    .io_count(mimoQ_io_count)
  );
  Computation compUnit_0 ( // @[programmableCache.scala 177:27]
    .clock(compUnit_0_clock),
    .reset(compUnit_0_reset),
    .io_instruction_valid(compUnit_0_io_instruction_valid),
    .io_instruction_bits(compUnit_0_io_instruction_bits),
    .io_clear(compUnit_0_io_clear),
    .io_op1_valid(compUnit_0_io_op1_valid),
    .io_op1_bits(compUnit_0_io_op1_bits),
    .io_op2_valid(compUnit_0_io_op2_valid),
    .io_op2_bits(compUnit_0_io_op2_bits),
    .io_pc(compUnit_0_io_pc),
    .io_reg_file_0(compUnit_0_io_reg_file_0),
    .io_reg_file_1(compUnit_0_io_reg_file_1),
    .io_reg_file_2(compUnit_0_io_reg_file_2),
    .io_reg_file_3(compUnit_0_io_reg_file_3)
  );
  Computation compUnit_1 ( // @[programmableCache.scala 177:27]
    .clock(compUnit_1_clock),
    .reset(compUnit_1_reset),
    .io_instruction_valid(compUnit_1_io_instruction_valid),
    .io_instruction_bits(compUnit_1_io_instruction_bits),
    .io_clear(compUnit_1_io_clear),
    .io_op1_valid(compUnit_1_io_op1_valid),
    .io_op1_bits(compUnit_1_io_op1_bits),
    .io_op2_valid(compUnit_1_io_op2_valid),
    .io_op2_bits(compUnit_1_io_op2_bits),
    .io_pc(compUnit_1_io_pc),
    .io_reg_file_0(compUnit_1_io_reg_file_0),
    .io_reg_file_1(compUnit_1_io_reg_file_1),
    .io_reg_file_2(compUnit_1_io_reg_file_2),
    .io_reg_file_3(compUnit_1_io_reg_file_3)
  );
  Computation compUnit_2 ( // @[programmableCache.scala 177:27]
    .clock(compUnit_2_clock),
    .reset(compUnit_2_reset),
    .io_instruction_valid(compUnit_2_io_instruction_valid),
    .io_instruction_bits(compUnit_2_io_instruction_bits),
    .io_clear(compUnit_2_io_clear),
    .io_op1_valid(compUnit_2_io_op1_valid),
    .io_op1_bits(compUnit_2_io_op1_bits),
    .io_op2_valid(compUnit_2_io_op2_valid),
    .io_op2_bits(compUnit_2_io_op2_bits),
    .io_pc(compUnit_2_io_pc),
    .io_reg_file_0(compUnit_2_io_reg_file_0),
    .io_reg_file_1(compUnit_2_io_reg_file_1),
    .io_reg_file_2(compUnit_2_io_reg_file_2),
    .io_reg_file_3(compUnit_2_io_reg_file_3)
  );
  Computation compUnit_3 ( // @[programmableCache.scala 177:27]
    .clock(compUnit_3_clock),
    .reset(compUnit_3_reset),
    .io_instruction_valid(compUnit_3_io_instruction_valid),
    .io_instruction_bits(compUnit_3_io_instruction_bits),
    .io_clear(compUnit_3_io_clear),
    .io_op1_valid(compUnit_3_io_op1_valid),
    .io_op1_bits(compUnit_3_io_op1_bits),
    .io_op2_valid(compUnit_3_io_op2_valid),
    .io_op2_bits(compUnit_3_io_op2_bits),
    .io_pc(compUnit_3_io_pc),
    .io_reg_file_0(compUnit_3_io_reg_file_0),
    .io_reg_file_1(compUnit_3_io_reg_file_1),
    .io_reg_file_2(compUnit_3_io_reg_file_2),
    .io_reg_file_3(compUnit_3_io_reg_file_3)
  );
  Computation compUnit_4 ( // @[programmableCache.scala 177:27]
    .clock(compUnit_4_clock),
    .reset(compUnit_4_reset),
    .io_instruction_valid(compUnit_4_io_instruction_valid),
    .io_instruction_bits(compUnit_4_io_instruction_bits),
    .io_clear(compUnit_4_io_clear),
    .io_op1_valid(compUnit_4_io_op1_valid),
    .io_op1_bits(compUnit_4_io_op1_bits),
    .io_op2_valid(compUnit_4_io_op2_valid),
    .io_op2_bits(compUnit_4_io_op2_bits),
    .io_pc(compUnit_4_io_pc),
    .io_reg_file_0(compUnit_4_io_reg_file_0),
    .io_reg_file_1(compUnit_4_io_reg_file_1),
    .io_reg_file_2(compUnit_4_io_reg_file_2),
    .io_reg_file_3(compUnit_4_io_reg_file_3)
  );
  Computation compUnit_5 ( // @[programmableCache.scala 177:27]
    .clock(compUnit_5_clock),
    .reset(compUnit_5_reset),
    .io_instruction_valid(compUnit_5_io_instruction_valid),
    .io_instruction_bits(compUnit_5_io_instruction_bits),
    .io_clear(compUnit_5_io_clear),
    .io_op1_valid(compUnit_5_io_op1_valid),
    .io_op1_bits(compUnit_5_io_op1_bits),
    .io_op2_valid(compUnit_5_io_op2_valid),
    .io_op2_bits(compUnit_5_io_op2_bits),
    .io_pc(compUnit_5_io_pc),
    .io_reg_file_0(compUnit_5_io_reg_file_0),
    .io_reg_file_1(compUnit_5_io_reg_file_1),
    .io_reg_file_2(compUnit_5_io_reg_file_2),
    .io_reg_file_3(compUnit_5_io_reg_file_3)
  );
  Computation compUnit_6 ( // @[programmableCache.scala 177:27]
    .clock(compUnit_6_clock),
    .reset(compUnit_6_reset),
    .io_instruction_valid(compUnit_6_io_instruction_valid),
    .io_instruction_bits(compUnit_6_io_instruction_bits),
    .io_clear(compUnit_6_io_clear),
    .io_op1_valid(compUnit_6_io_op1_valid),
    .io_op1_bits(compUnit_6_io_op1_bits),
    .io_op2_valid(compUnit_6_io_op2_valid),
    .io_op2_bits(compUnit_6_io_op2_bits),
    .io_pc(compUnit_6_io_pc),
    .io_reg_file_0(compUnit_6_io_reg_file_0),
    .io_reg_file_1(compUnit_6_io_reg_file_1),
    .io_reg_file_2(compUnit_6_io_reg_file_2),
    .io_reg_file_3(compUnit_6_io_reg_file_3)
  );
  Computation compUnit_7 ( // @[programmableCache.scala 177:27]
    .clock(compUnit_7_clock),
    .reset(compUnit_7_reset),
    .io_instruction_valid(compUnit_7_io_instruction_valid),
    .io_instruction_bits(compUnit_7_io_instruction_bits),
    .io_clear(compUnit_7_io_clear),
    .io_op1_valid(compUnit_7_io_op1_valid),
    .io_op1_bits(compUnit_7_io_op1_bits),
    .io_op2_valid(compUnit_7_io_op2_valid),
    .io_op2_bits(compUnit_7_io_op2_bits),
    .io_pc(compUnit_7_io_pc),
    .io_reg_file_0(compUnit_7_io_reg_file_0),
    .io_reg_file_1(compUnit_7_io_reg_file_1),
    .io_reg_file_2(compUnit_7_io_reg_file_2),
    .io_reg_file_3(compUnit_7_io_reg_file_3)
  );
  Mux3 compUnitInput1_0 ( // @[programmableCache.scala 182:30]
    .io_in_hardCoded(compUnitInput1_0_io_in_hardCoded),
    .io_in_data(compUnitInput1_0_io_in_data),
    .io_in_tbe(compUnitInput1_0_io_in_tbe),
    .io_in_select(compUnitInput1_0_io_in_select),
    .io_out_valid(compUnitInput1_0_io_out_valid),
    .io_out_bits(compUnitInput1_0_io_out_bits)
  );
  Mux3 compUnitInput1_1 ( // @[programmableCache.scala 182:30]
    .io_in_hardCoded(compUnitInput1_1_io_in_hardCoded),
    .io_in_data(compUnitInput1_1_io_in_data),
    .io_in_tbe(compUnitInput1_1_io_in_tbe),
    .io_in_select(compUnitInput1_1_io_in_select),
    .io_out_valid(compUnitInput1_1_io_out_valid),
    .io_out_bits(compUnitInput1_1_io_out_bits)
  );
  Mux3 compUnitInput1_2 ( // @[programmableCache.scala 182:30]
    .io_in_hardCoded(compUnitInput1_2_io_in_hardCoded),
    .io_in_data(compUnitInput1_2_io_in_data),
    .io_in_tbe(compUnitInput1_2_io_in_tbe),
    .io_in_select(compUnitInput1_2_io_in_select),
    .io_out_valid(compUnitInput1_2_io_out_valid),
    .io_out_bits(compUnitInput1_2_io_out_bits)
  );
  Mux3 compUnitInput1_3 ( // @[programmableCache.scala 182:30]
    .io_in_hardCoded(compUnitInput1_3_io_in_hardCoded),
    .io_in_data(compUnitInput1_3_io_in_data),
    .io_in_tbe(compUnitInput1_3_io_in_tbe),
    .io_in_select(compUnitInput1_3_io_in_select),
    .io_out_valid(compUnitInput1_3_io_out_valid),
    .io_out_bits(compUnitInput1_3_io_out_bits)
  );
  Mux3 compUnitInput1_4 ( // @[programmableCache.scala 182:30]
    .io_in_hardCoded(compUnitInput1_4_io_in_hardCoded),
    .io_in_data(compUnitInput1_4_io_in_data),
    .io_in_tbe(compUnitInput1_4_io_in_tbe),
    .io_in_select(compUnitInput1_4_io_in_select),
    .io_out_valid(compUnitInput1_4_io_out_valid),
    .io_out_bits(compUnitInput1_4_io_out_bits)
  );
  Mux3 compUnitInput1_5 ( // @[programmableCache.scala 182:30]
    .io_in_hardCoded(compUnitInput1_5_io_in_hardCoded),
    .io_in_data(compUnitInput1_5_io_in_data),
    .io_in_tbe(compUnitInput1_5_io_in_tbe),
    .io_in_select(compUnitInput1_5_io_in_select),
    .io_out_valid(compUnitInput1_5_io_out_valid),
    .io_out_bits(compUnitInput1_5_io_out_bits)
  );
  Mux3 compUnitInput1_6 ( // @[programmableCache.scala 182:30]
    .io_in_hardCoded(compUnitInput1_6_io_in_hardCoded),
    .io_in_data(compUnitInput1_6_io_in_data),
    .io_in_tbe(compUnitInput1_6_io_in_tbe),
    .io_in_select(compUnitInput1_6_io_in_select),
    .io_out_valid(compUnitInput1_6_io_out_valid),
    .io_out_bits(compUnitInput1_6_io_out_bits)
  );
  Mux3 compUnitInput1_7 ( // @[programmableCache.scala 182:30]
    .io_in_hardCoded(compUnitInput1_7_io_in_hardCoded),
    .io_in_data(compUnitInput1_7_io_in_data),
    .io_in_tbe(compUnitInput1_7_io_in_tbe),
    .io_in_select(compUnitInput1_7_io_in_select),
    .io_out_valid(compUnitInput1_7_io_out_valid),
    .io_out_bits(compUnitInput1_7_io_out_bits)
  );
  Mux3 compUnitInput2_0 ( // @[programmableCache.scala 188:30]
    .io_in_hardCoded(compUnitInput2_0_io_in_hardCoded),
    .io_in_data(compUnitInput2_0_io_in_data),
    .io_in_tbe(compUnitInput2_0_io_in_tbe),
    .io_in_select(compUnitInput2_0_io_in_select),
    .io_out_valid(compUnitInput2_0_io_out_valid),
    .io_out_bits(compUnitInput2_0_io_out_bits)
  );
  Mux3 compUnitInput2_1 ( // @[programmableCache.scala 188:30]
    .io_in_hardCoded(compUnitInput2_1_io_in_hardCoded),
    .io_in_data(compUnitInput2_1_io_in_data),
    .io_in_tbe(compUnitInput2_1_io_in_tbe),
    .io_in_select(compUnitInput2_1_io_in_select),
    .io_out_valid(compUnitInput2_1_io_out_valid),
    .io_out_bits(compUnitInput2_1_io_out_bits)
  );
  Mux3 compUnitInput2_2 ( // @[programmableCache.scala 188:30]
    .io_in_hardCoded(compUnitInput2_2_io_in_hardCoded),
    .io_in_data(compUnitInput2_2_io_in_data),
    .io_in_tbe(compUnitInput2_2_io_in_tbe),
    .io_in_select(compUnitInput2_2_io_in_select),
    .io_out_valid(compUnitInput2_2_io_out_valid),
    .io_out_bits(compUnitInput2_2_io_out_bits)
  );
  Mux3 compUnitInput2_3 ( // @[programmableCache.scala 188:30]
    .io_in_hardCoded(compUnitInput2_3_io_in_hardCoded),
    .io_in_data(compUnitInput2_3_io_in_data),
    .io_in_tbe(compUnitInput2_3_io_in_tbe),
    .io_in_select(compUnitInput2_3_io_in_select),
    .io_out_valid(compUnitInput2_3_io_out_valid),
    .io_out_bits(compUnitInput2_3_io_out_bits)
  );
  Mux3 compUnitInput2_4 ( // @[programmableCache.scala 188:30]
    .io_in_hardCoded(compUnitInput2_4_io_in_hardCoded),
    .io_in_data(compUnitInput2_4_io_in_data),
    .io_in_tbe(compUnitInput2_4_io_in_tbe),
    .io_in_select(compUnitInput2_4_io_in_select),
    .io_out_valid(compUnitInput2_4_io_out_valid),
    .io_out_bits(compUnitInput2_4_io_out_bits)
  );
  Mux3 compUnitInput2_5 ( // @[programmableCache.scala 188:30]
    .io_in_hardCoded(compUnitInput2_5_io_in_hardCoded),
    .io_in_data(compUnitInput2_5_io_in_data),
    .io_in_tbe(compUnitInput2_5_io_in_tbe),
    .io_in_select(compUnitInput2_5_io_in_select),
    .io_out_valid(compUnitInput2_5_io_out_valid),
    .io_out_bits(compUnitInput2_5_io_out_bits)
  );
  Mux3 compUnitInput2_6 ( // @[programmableCache.scala 188:30]
    .io_in_hardCoded(compUnitInput2_6_io_in_hardCoded),
    .io_in_data(compUnitInput2_6_io_in_data),
    .io_in_tbe(compUnitInput2_6_io_in_tbe),
    .io_in_select(compUnitInput2_6_io_in_select),
    .io_out_valid(compUnitInput2_6_io_out_valid),
    .io_out_bits(compUnitInput2_6_io_out_bits)
  );
  Mux3 compUnitInput2_7 ( // @[programmableCache.scala 188:30]
    .io_in_hardCoded(compUnitInput2_7_io_in_hardCoded),
    .io_in_data(compUnitInput2_7_io_in_data),
    .io_in_tbe(compUnitInput2_7_io_in_tbe),
    .io_in_select(compUnitInput2_7_io_in_select),
    .io_out_valid(compUnitInput2_7_io_out_valid),
    .io_out_bits(compUnitInput2_7_io_out_bits)
  );
  assign io_in_cpu_ready = _T_141 & _T_161; // @[programmableCache.scala 240:37 programmableCache.scala 280:28]
  assign io_in_memCtrl_ready = _T_141 & _T_158; // @[programmableCache.scala 241:41 programmableCache.scala 279:28]
  assign io_in_otherNodes_ready = _T_141 & _T_164; // @[programmableCache.scala 239:44 programmableCache.scala 281:28]
  assign io_out_req_valid = outReqArbiter_io_out_valid; // @[programmableCache.scala 499:22]
  assign io_out_req_bits_req_addr = outReqArbiter_io_out_bits_req_addr; // @[programmableCache.scala 497:30]
  assign io_out_req_bits_req_inst = outReqArbiter_io_out_bits_req_inst; // @[programmableCache.scala 495:30]
  assign io_out_req_bits_req_data = outReqArbiter_io_out_bits_req_data; // @[programmableCache.scala 496:30]
  assign io_out_resp_valid = outRespArbiter_io_out_valid; // @[programmableCache.scala 525:27]
  assign io_out_resp_bits_addr = outRespArbiter_io_out_bits_addr; // @[programmableCache.scala 524:27]
  assign _T_814_0 = _T_159;
  assign _T_808_0 = _T_141;
  assign _T_819_0 = probeStart;
  assign hitLD_0 = hitLD;
  assign missLD_0 = missLD;
  assign _T_811_0 = _T_162;
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_cpu_0_req_valid = actionReg_0_io_deq_ready & actionReg_0_io_deq_valid; // @[programmableCache.scala 460:35]
  assign cache_io_cpu_0_req_bits_addr = actionReg_0_io_deq_bits_addr; // @[programmableCache.scala 459:39]
  assign cache_io_cpu_0_req_bits_command = isCacheAction_0 ? actionReg_0_io_deq_bits_action_signals : 28'h0; // @[programmableCache.scala 458:42]
  assign cache_io_cpu_0_req_bits_way = actionReg_0_io_deq_bits_way; // @[programmableCache.scala 457:38]
  assign cache_io_cpu_0_req_bits_replaceWay = actionReg_0_io_deq_bits_replaceWay; // @[programmableCache.scala 462:45]
  assign cache_io_cpu_1_req_valid = actionReg_1_io_deq_ready & actionReg_1_io_deq_valid; // @[programmableCache.scala 460:35]
  assign cache_io_cpu_1_req_bits_addr = actionReg_1_io_deq_bits_addr; // @[programmableCache.scala 459:39]
  assign cache_io_cpu_1_req_bits_command = isCacheAction_1 ? actionReg_1_io_deq_bits_action_signals : 28'h0; // @[programmableCache.scala 458:42]
  assign cache_io_cpu_1_req_bits_way = actionReg_1_io_deq_bits_way; // @[programmableCache.scala 457:38]
  assign cache_io_cpu_1_req_bits_replaceWay = actionReg_1_io_deq_bits_replaceWay; // @[programmableCache.scala 462:45]
  assign cache_io_cpu_2_req_valid = actionReg_2_io_deq_ready & actionReg_2_io_deq_valid; // @[programmableCache.scala 460:35]
  assign cache_io_cpu_2_req_bits_addr = actionReg_2_io_deq_bits_addr; // @[programmableCache.scala 459:39]
  assign cache_io_cpu_2_req_bits_command = isCacheAction_2 ? actionReg_2_io_deq_bits_action_signals : 28'h0; // @[programmableCache.scala 458:42]
  assign cache_io_cpu_2_req_bits_way = actionReg_2_io_deq_bits_way; // @[programmableCache.scala 457:38]
  assign cache_io_cpu_2_req_bits_replaceWay = actionReg_2_io_deq_bits_replaceWay; // @[programmableCache.scala 462:45]
  assign cache_io_cpu_3_req_valid = actionReg_3_io_deq_ready & actionReg_3_io_deq_valid; // @[programmableCache.scala 460:35]
  assign cache_io_cpu_3_req_bits_addr = actionReg_3_io_deq_bits_addr; // @[programmableCache.scala 459:39]
  assign cache_io_cpu_3_req_bits_command = isCacheAction_3 ? actionReg_3_io_deq_bits_action_signals : 28'h0; // @[programmableCache.scala 458:42]
  assign cache_io_cpu_3_req_bits_way = actionReg_3_io_deq_bits_way; // @[programmableCache.scala 457:38]
  assign cache_io_cpu_3_req_bits_replaceWay = actionReg_3_io_deq_bits_replaceWay; // @[programmableCache.scala 462:45]
  assign cache_io_cpu_4_req_valid = actionReg_4_io_deq_ready & actionReg_4_io_deq_valid; // @[programmableCache.scala 460:35]
  assign cache_io_cpu_4_req_bits_addr = actionReg_4_io_deq_bits_addr; // @[programmableCache.scala 459:39]
  assign cache_io_cpu_4_req_bits_command = isCacheAction_4 ? actionReg_4_io_deq_bits_action_signals : 28'h0; // @[programmableCache.scala 458:42]
  assign cache_io_cpu_4_req_bits_way = actionReg_4_io_deq_bits_way; // @[programmableCache.scala 457:38]
  assign cache_io_cpu_4_req_bits_replaceWay = actionReg_4_io_deq_bits_replaceWay; // @[programmableCache.scala 462:45]
  assign cache_io_cpu_5_req_valid = actionReg_5_io_deq_ready & actionReg_5_io_deq_valid; // @[programmableCache.scala 460:35]
  assign cache_io_cpu_5_req_bits_addr = actionReg_5_io_deq_bits_addr; // @[programmableCache.scala 459:39]
  assign cache_io_cpu_5_req_bits_command = isCacheAction_5 ? actionReg_5_io_deq_bits_action_signals : 28'h0; // @[programmableCache.scala 458:42]
  assign cache_io_cpu_5_req_bits_way = actionReg_5_io_deq_bits_way; // @[programmableCache.scala 457:38]
  assign cache_io_cpu_5_req_bits_replaceWay = actionReg_5_io_deq_bits_replaceWay; // @[programmableCache.scala 462:45]
  assign cache_io_cpu_6_req_valid = actionReg_6_io_deq_ready & actionReg_6_io_deq_valid; // @[programmableCache.scala 460:35]
  assign cache_io_cpu_6_req_bits_addr = actionReg_6_io_deq_bits_addr; // @[programmableCache.scala 459:39]
  assign cache_io_cpu_6_req_bits_command = isCacheAction_6 ? actionReg_6_io_deq_bits_action_signals : 28'h0; // @[programmableCache.scala 458:42]
  assign cache_io_cpu_6_req_bits_way = actionReg_6_io_deq_bits_way; // @[programmableCache.scala 457:38]
  assign cache_io_cpu_6_req_bits_replaceWay = actionReg_6_io_deq_bits_replaceWay; // @[programmableCache.scala 462:45]
  assign cache_io_cpu_7_req_valid = actionReg_7_io_deq_ready & actionReg_7_io_deq_valid; // @[programmableCache.scala 460:35]
  assign cache_io_cpu_7_req_bits_addr = actionReg_7_io_deq_bits_addr; // @[programmableCache.scala 459:39]
  assign cache_io_cpu_7_req_bits_data = actionReg_7_io_deq_bits_data; // @[programmableCache.scala 461:39]
  assign cache_io_cpu_7_req_bits_command = isCacheAction_7 ? actionReg_7_io_deq_bits_action_signals : 28'h0; // @[programmableCache.scala 458:42]
  assign cache_io_cpu_7_req_bits_way = actionReg_7_io_deq_bits_way; // @[programmableCache.scala 457:38]
  assign cache_io_cpu_7_req_bits_replaceWay = actionReg_7_io_deq_bits_replaceWay; // @[programmableCache.scala 462:45]
  assign cache_io_probe_req_valid = _T_141 & _T_142; // @[programmableCache.scala 468:30]
  assign cache_io_probe_req_bits_addr = probeStart ? instruction_bits_addr : 32'h0; // @[programmableCache.scala 466:34]
  assign cache_io_probe_req_bits_command = probeStart ? 28'hb : 28'h0; // @[programmableCache.scala 465:37]
  assign cache_io_bipassLD_in_valid = mimoQ_io_deq_valid & _T_741; // @[programmableCache.scala 471:32]
  assign cache_io_bipassLD_in_bits_addr = mimoQ_io_deq_bits_0_addr; // @[programmableCache.scala 472:37]
  assign cache_io_bipassLD_in_bits_way = {{1'd0}, mimoQ_io_deq_bits_0_way}; // @[programmableCache.scala 473:35]
  assign tbe_clock = clock;
  assign tbe_reset = reset;
  assign tbe_io_write_0_valid = isTBEAction_0 | isStateAction_0; // @[programmableCache.scala 309:31]
  assign tbe_io_write_0_bits_addr = {{32'd0}, actionReg_0_io_deq_bits_addr}; // @[programmableCache.scala 306:35]
  assign tbe_io_write_0_bits_command = isStateAction_0 ? 2'h3 : tbeAction_0; // @[programmableCache.scala 305:38]
  assign tbe_io_write_0_bits_mask = isStateAction_0 | maskField_0; // @[programmableCache.scala 308:35]
  assign tbe_io_write_0_bits_inputTBE_state_state = isStateAction_0 ? tbeAction_0 : 2'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_0_bits_inputTBE_way = {{1'd0}, actionReg_0_io_deq_bits_way}; // @[programmableCache.scala 307:39]
  assign tbe_io_write_0_bits_inputTBE_fields_0 = _T_185 ? tbeFieldUpdateSrc_0 : 32'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_1_valid = isTBEAction_1 | isStateAction_1; // @[programmableCache.scala 309:31]
  assign tbe_io_write_1_bits_addr = {{32'd0}, actionReg_1_io_deq_bits_addr}; // @[programmableCache.scala 306:35]
  assign tbe_io_write_1_bits_command = isStateAction_1 ? 2'h3 : tbeAction_1; // @[programmableCache.scala 305:38]
  assign tbe_io_write_1_bits_mask = isStateAction_1 | maskField_1; // @[programmableCache.scala 308:35]
  assign tbe_io_write_1_bits_inputTBE_state_state = isStateAction_1 ? tbeAction_1 : 2'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_1_bits_inputTBE_way = {{1'd0}, actionReg_1_io_deq_bits_way}; // @[programmableCache.scala 307:39]
  assign tbe_io_write_1_bits_inputTBE_fields_0 = _T_191 ? tbeFieldUpdateSrc_1 : 32'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_2_valid = isTBEAction_2 | isStateAction_2; // @[programmableCache.scala 309:31]
  assign tbe_io_write_2_bits_addr = {{32'd0}, actionReg_2_io_deq_bits_addr}; // @[programmableCache.scala 306:35]
  assign tbe_io_write_2_bits_command = isStateAction_2 ? 2'h3 : tbeAction_2; // @[programmableCache.scala 305:38]
  assign tbe_io_write_2_bits_mask = isStateAction_2 | maskField_2; // @[programmableCache.scala 308:35]
  assign tbe_io_write_2_bits_inputTBE_state_state = isStateAction_2 ? tbeAction_2 : 2'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_2_bits_inputTBE_way = {{1'd0}, actionReg_2_io_deq_bits_way}; // @[programmableCache.scala 307:39]
  assign tbe_io_write_2_bits_inputTBE_fields_0 = _T_197 ? tbeFieldUpdateSrc_2 : 32'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_3_valid = isTBEAction_3 | isStateAction_3; // @[programmableCache.scala 309:31]
  assign tbe_io_write_3_bits_addr = {{32'd0}, actionReg_3_io_deq_bits_addr}; // @[programmableCache.scala 306:35]
  assign tbe_io_write_3_bits_command = isStateAction_3 ? 2'h3 : tbeAction_3; // @[programmableCache.scala 305:38]
  assign tbe_io_write_3_bits_mask = isStateAction_3 | maskField_3; // @[programmableCache.scala 308:35]
  assign tbe_io_write_3_bits_inputTBE_state_state = isStateAction_3 ? tbeAction_3 : 2'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_3_bits_inputTBE_way = {{1'd0}, actionReg_3_io_deq_bits_way}; // @[programmableCache.scala 307:39]
  assign tbe_io_write_3_bits_inputTBE_fields_0 = _T_203 ? tbeFieldUpdateSrc_3 : 32'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_4_valid = isTBEAction_4 | isStateAction_4; // @[programmableCache.scala 309:31]
  assign tbe_io_write_4_bits_addr = {{32'd0}, actionReg_4_io_deq_bits_addr}; // @[programmableCache.scala 306:35]
  assign tbe_io_write_4_bits_command = isStateAction_4 ? 2'h3 : tbeAction_4; // @[programmableCache.scala 305:38]
  assign tbe_io_write_4_bits_mask = isStateAction_4 | maskField_4; // @[programmableCache.scala 308:35]
  assign tbe_io_write_4_bits_inputTBE_state_state = isStateAction_4 ? tbeAction_4 : 2'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_4_bits_inputTBE_way = {{1'd0}, actionReg_4_io_deq_bits_way}; // @[programmableCache.scala 307:39]
  assign tbe_io_write_4_bits_inputTBE_fields_0 = _T_209 ? tbeFieldUpdateSrc_4 : 32'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_5_valid = isTBEAction_5 | isStateAction_5; // @[programmableCache.scala 309:31]
  assign tbe_io_write_5_bits_addr = {{32'd0}, actionReg_5_io_deq_bits_addr}; // @[programmableCache.scala 306:35]
  assign tbe_io_write_5_bits_command = isStateAction_5 ? 2'h3 : tbeAction_5; // @[programmableCache.scala 305:38]
  assign tbe_io_write_5_bits_mask = isStateAction_5 | maskField_5; // @[programmableCache.scala 308:35]
  assign tbe_io_write_5_bits_inputTBE_state_state = isStateAction_5 ? tbeAction_5 : 2'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_5_bits_inputTBE_way = {{1'd0}, actionReg_5_io_deq_bits_way}; // @[programmableCache.scala 307:39]
  assign tbe_io_write_5_bits_inputTBE_fields_0 = _T_215 ? tbeFieldUpdateSrc_5 : 32'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_6_valid = isTBEAction_6 | isStateAction_6; // @[programmableCache.scala 309:31]
  assign tbe_io_write_6_bits_addr = {{32'd0}, actionReg_6_io_deq_bits_addr}; // @[programmableCache.scala 306:35]
  assign tbe_io_write_6_bits_command = isStateAction_6 ? 2'h3 : tbeAction_6; // @[programmableCache.scala 305:38]
  assign tbe_io_write_6_bits_mask = isStateAction_6 | maskField_6; // @[programmableCache.scala 308:35]
  assign tbe_io_write_6_bits_inputTBE_state_state = isStateAction_6 ? tbeAction_6 : 2'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_6_bits_inputTBE_way = {{1'd0}, actionReg_6_io_deq_bits_way}; // @[programmableCache.scala 307:39]
  assign tbe_io_write_6_bits_inputTBE_fields_0 = _T_221 ? tbeFieldUpdateSrc_6 : 32'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_7_valid = isTBEAction_7 | isStateAction_7; // @[programmableCache.scala 309:31]
  assign tbe_io_write_7_bits_addr = {{32'd0}, actionReg_7_io_deq_bits_addr}; // @[programmableCache.scala 306:35]
  assign tbe_io_write_7_bits_command = isStateAction_7 ? 2'h3 : tbeAction_7; // @[programmableCache.scala 305:38]
  assign tbe_io_write_7_bits_mask = isStateAction_7 | maskField_7; // @[programmableCache.scala 308:35]
  assign tbe_io_write_7_bits_inputTBE_state_state = isStateAction_7 ? tbeAction_7 : 2'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_7_bits_inputTBE_way = {{1'd0}, actionReg_7_io_deq_bits_way}; // @[programmableCache.scala 307:39]
  assign tbe_io_write_7_bits_inputTBE_fields_0 = _T_227 ? tbeFieldUpdateSrc_7 : 32'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_read_valid = inputArbiter_io_out_valid; // @[programmableCache.scala 297:23]
  assign tbe_io_read_bits_addr = {{32'd0}, inputArbiter_io_out_bits_addr}; // @[programmableCache.scala 298:27]
  assign lockMem_clock = clock;
  assign lockMem_reset = reset;
  assign lockMem_io_lock_in_valid = instruction_ready & instruction_valid; // @[programmableCache.scala 320:35]
  assign lockMem_io_lock_in_bits_addr = inputArbiter_io_out_bits_addr; // @[programmableCache.scala 319:35]
  assign lockMem_io_probe_in_valid = inputArbiter_io_out_valid; // @[programmableCache.scala 315:35]
  assign lockMem_io_probe_in_bits_addr = inputArbiter_io_out_bits_addr; // @[programmableCache.scala 314:35]
  assign lockMem_io_unLock_0_in_valid = _T_280 & actionReg_0_io_deq_valid; // @[programmableCache.scala 328:39]
  assign lockMem_io_unLock_0_in_bits_addr = actionReg_0_io_deq_bits_addr; // @[programmableCache.scala 326:43]
  assign lockMem_io_unLock_1_in_valid = _T_337 & actionReg_1_io_deq_valid; // @[programmableCache.scala 328:39]
  assign lockMem_io_unLock_1_in_bits_addr = actionReg_1_io_deq_bits_addr; // @[programmableCache.scala 326:43]
  assign lockMem_io_unLock_2_in_valid = _T_394 & actionReg_2_io_deq_valid; // @[programmableCache.scala 328:39]
  assign lockMem_io_unLock_2_in_bits_addr = actionReg_2_io_deq_bits_addr; // @[programmableCache.scala 326:43]
  assign lockMem_io_unLock_3_in_valid = _T_451 & actionReg_3_io_deq_valid; // @[programmableCache.scala 328:39]
  assign lockMem_io_unLock_3_in_bits_addr = actionReg_3_io_deq_bits_addr; // @[programmableCache.scala 326:43]
  assign lockMem_io_unLock_4_in_valid = _T_508 & actionReg_4_io_deq_valid; // @[programmableCache.scala 328:39]
  assign lockMem_io_unLock_4_in_bits_addr = actionReg_4_io_deq_bits_addr; // @[programmableCache.scala 326:43]
  assign lockMem_io_unLock_5_in_valid = _T_565 & actionReg_5_io_deq_valid; // @[programmableCache.scala 328:39]
  assign lockMem_io_unLock_5_in_bits_addr = actionReg_5_io_deq_bits_addr; // @[programmableCache.scala 326:43]
  assign lockMem_io_unLock_6_in_valid = _T_622 & actionReg_6_io_deq_valid; // @[programmableCache.scala 328:39]
  assign lockMem_io_unLock_6_in_bits_addr = actionReg_6_io_deq_bits_addr; // @[programmableCache.scala 326:43]
  assign lockMem_io_unLock_7_in_valid = _T_679 & actionReg_7_io_deq_valid; // @[programmableCache.scala 328:39]
  assign lockMem_io_unLock_7_in_bits_addr = actionReg_7_io_deq_bits_addr; // @[programmableCache.scala 326:43]
  assign stateMem_clock = clock;
  assign stateMem_reset = reset;
  assign stateMem_io_in_0_valid = _T_280 & actionReg_0_io_deq_valid; // @[programmableCache.scala 338:33]
  assign stateMem_io_in_0_bits_state_state = isStateAction_0 ? tbeAction_0 : 2'h0; // @[programmableCache.scala 336:38]
  assign stateMem_io_in_0_bits_addr = actionReg_0_io_deq_bits_addr; // @[programmableCache.scala 335:37]
  assign stateMem_io_in_0_bits_way = actionReg_0_io_deq_bits_way; // @[programmableCache.scala 337:36]
  assign stateMem_io_in_1_valid = _T_337 & actionReg_1_io_deq_valid; // @[programmableCache.scala 338:33]
  assign stateMem_io_in_1_bits_state_state = isStateAction_1 ? tbeAction_1 : 2'h0; // @[programmableCache.scala 336:38]
  assign stateMem_io_in_1_bits_addr = actionReg_1_io_deq_bits_addr; // @[programmableCache.scala 335:37]
  assign stateMem_io_in_1_bits_way = actionReg_1_io_deq_bits_way; // @[programmableCache.scala 337:36]
  assign stateMem_io_in_2_valid = _T_394 & actionReg_2_io_deq_valid; // @[programmableCache.scala 338:33]
  assign stateMem_io_in_2_bits_state_state = isStateAction_2 ? tbeAction_2 : 2'h0; // @[programmableCache.scala 336:38]
  assign stateMem_io_in_2_bits_addr = actionReg_2_io_deq_bits_addr; // @[programmableCache.scala 335:37]
  assign stateMem_io_in_2_bits_way = actionReg_2_io_deq_bits_way; // @[programmableCache.scala 337:36]
  assign stateMem_io_in_3_valid = _T_451 & actionReg_3_io_deq_valid; // @[programmableCache.scala 338:33]
  assign stateMem_io_in_3_bits_state_state = isStateAction_3 ? tbeAction_3 : 2'h0; // @[programmableCache.scala 336:38]
  assign stateMem_io_in_3_bits_addr = actionReg_3_io_deq_bits_addr; // @[programmableCache.scala 335:37]
  assign stateMem_io_in_3_bits_way = actionReg_3_io_deq_bits_way; // @[programmableCache.scala 337:36]
  assign stateMem_io_in_4_valid = _T_508 & actionReg_4_io_deq_valid; // @[programmableCache.scala 338:33]
  assign stateMem_io_in_4_bits_state_state = isStateAction_4 ? tbeAction_4 : 2'h0; // @[programmableCache.scala 336:38]
  assign stateMem_io_in_4_bits_addr = actionReg_4_io_deq_bits_addr; // @[programmableCache.scala 335:37]
  assign stateMem_io_in_4_bits_way = actionReg_4_io_deq_bits_way; // @[programmableCache.scala 337:36]
  assign stateMem_io_in_5_valid = _T_565 & actionReg_5_io_deq_valid; // @[programmableCache.scala 338:33]
  assign stateMem_io_in_5_bits_state_state = isStateAction_5 ? tbeAction_5 : 2'h0; // @[programmableCache.scala 336:38]
  assign stateMem_io_in_5_bits_addr = actionReg_5_io_deq_bits_addr; // @[programmableCache.scala 335:37]
  assign stateMem_io_in_5_bits_way = actionReg_5_io_deq_bits_way; // @[programmableCache.scala 337:36]
  assign stateMem_io_in_6_valid = _T_622 & actionReg_6_io_deq_valid; // @[programmableCache.scala 338:33]
  assign stateMem_io_in_6_bits_state_state = isStateAction_6 ? tbeAction_6 : 2'h0; // @[programmableCache.scala 336:38]
  assign stateMem_io_in_6_bits_addr = actionReg_6_io_deq_bits_addr; // @[programmableCache.scala 335:37]
  assign stateMem_io_in_6_bits_way = actionReg_6_io_deq_bits_way; // @[programmableCache.scala 337:36]
  assign stateMem_io_in_7_valid = _T_679 & actionReg_7_io_deq_valid; // @[programmableCache.scala 338:33]
  assign stateMem_io_in_7_bits_state_state = isStateAction_7 ? tbeAction_7 : 2'h0; // @[programmableCache.scala 336:38]
  assign stateMem_io_in_7_bits_addr = actionReg_7_io_deq_bits_addr; // @[programmableCache.scala 335:37]
  assign stateMem_io_in_7_bits_way = actionReg_7_io_deq_bits_way; // @[programmableCache.scala 337:36]
  assign stateMem_io_in_8_valid = input__io_deq_ready & input__io_deq_valid; // @[programmableCache.scala 345:34]
  assign stateMem_io_in_8_bits_addr = input__io_deq_bits_inst_addr; // @[programmableCache.scala 342:38]
  assign stateMem_io_in_8_bits_way = probeWay_io_deq_bits; // @[programmableCache.scala 344:37]
  assign pc_clock = clock;
  assign pc_reset = reset;
  assign pc_io_write_valid = routineQueue_io_deq_ready & routineQueue_io_deq_valid; // @[programmableCache.scala 451:23]
  assign pc_io_write_bits_addr = inputToPC_addr; // @[programmableCache.scala 443:27]
  assign pc_io_write_bits_way = wayInputCache[1:0]; // @[programmableCache.scala 444:26]
  assign pc_io_write_bits_data = inputToPC_data; // @[programmableCache.scala 448:27]
  assign pc_io_write_bits_replaceWay = replaceWayInputCache[1:0]; // @[programmableCache.scala 446:33]
  assign pc_io_write_bits_tbeFields_0 = tbeFields_0; // @[programmableCache.scala 445:32]
  assign pc_io_write_bits_pc = routineQueue_io_deq_bits; // @[programmableCache.scala 447:25]
  assign pc_io_read_0_in_bits_data_way = _T_301[1:0]; // @[programmableCache.scala 398:40]
  assign pc_io_read_0_in_bits_data_pc = firstLineNextRoutine_0 ? pcWire_0_pc : _T_296; // @[programmableCache.scala 400:39]
  assign pc_io_read_0_in_bits_data_valid = ~firstLineNextRoutine_0; // @[programmableCache.scala 403:42]
  assign pc_io_read_1_in_bits_data_way = _T_358[1:0]; // @[programmableCache.scala 398:40]
  assign pc_io_read_1_in_bits_data_pc = firstLineNextRoutine_1 ? pcWire_1_pc : _T_353; // @[programmableCache.scala 400:39]
  assign pc_io_read_1_in_bits_data_valid = ~firstLineNextRoutine_1; // @[programmableCache.scala 403:42]
  assign pc_io_read_2_in_bits_data_way = _T_415[1:0]; // @[programmableCache.scala 398:40]
  assign pc_io_read_2_in_bits_data_pc = firstLineNextRoutine_2 ? pcWire_2_pc : _T_410; // @[programmableCache.scala 400:39]
  assign pc_io_read_2_in_bits_data_valid = ~firstLineNextRoutine_2; // @[programmableCache.scala 403:42]
  assign pc_io_read_3_in_bits_data_way = _T_472[1:0]; // @[programmableCache.scala 398:40]
  assign pc_io_read_3_in_bits_data_pc = firstLineNextRoutine_3 ? pcWire_3_pc : _T_467; // @[programmableCache.scala 400:39]
  assign pc_io_read_3_in_bits_data_valid = ~firstLineNextRoutine_3; // @[programmableCache.scala 403:42]
  assign pc_io_read_4_in_bits_data_way = _T_529[1:0]; // @[programmableCache.scala 398:40]
  assign pc_io_read_4_in_bits_data_pc = firstLineNextRoutine_4 ? pcWire_4_pc : _T_524; // @[programmableCache.scala 400:39]
  assign pc_io_read_4_in_bits_data_valid = ~firstLineNextRoutine_4; // @[programmableCache.scala 403:42]
  assign pc_io_read_5_in_bits_data_way = _T_586[1:0]; // @[programmableCache.scala 398:40]
  assign pc_io_read_5_in_bits_data_pc = firstLineNextRoutine_5 ? pcWire_5_pc : _T_581; // @[programmableCache.scala 400:39]
  assign pc_io_read_5_in_bits_data_valid = ~firstLineNextRoutine_5; // @[programmableCache.scala 403:42]
  assign pc_io_read_6_in_bits_data_way = _T_643[1:0]; // @[programmableCache.scala 398:40]
  assign pc_io_read_6_in_bits_data_pc = firstLineNextRoutine_6 ? pcWire_6_pc : _T_638; // @[programmableCache.scala 400:39]
  assign pc_io_read_6_in_bits_data_valid = ~firstLineNextRoutine_6; // @[programmableCache.scala 403:42]
  assign pc_io_read_7_in_bits_data_way = _T_700[1:0]; // @[programmableCache.scala 398:40]
  assign pc_io_read_7_in_bits_data_pc = firstLineNextRoutine_7 ? pcWire_7_pc : _T_695; // @[programmableCache.scala 400:39]
  assign pc_io_read_7_in_bits_data_valid = ~firstLineNextRoutine_7; // @[programmableCache.scala 403:42]
  assign inputArbiter_io_in_0_valid = io_in_memCtrl_valid; // @[programmableCache.scala 241:41]
  assign inputArbiter_io_in_0_bits_event = io_in_memCtrl_bits_event; // @[programmableCache.scala 241:41]
  assign inputArbiter_io_in_0_bits_addr = io_in_memCtrl_bits_addr; // @[programmableCache.scala 241:41]
  assign inputArbiter_io_in_0_bits_data = io_in_memCtrl_bits_data; // @[programmableCache.scala 241:41]
  assign inputArbiter_io_in_1_valid = feedbackOutQueue_io_deq_valid; // @[programmableCache.scala 242:42]
  assign inputArbiter_io_in_1_bits_event = feedbackOutQueue_io_deq_bits_event; // @[programmableCache.scala 242:42]
  assign inputArbiter_io_in_1_bits_addr = feedbackOutQueue_io_deq_bits_addr; // @[programmableCache.scala 242:42]
  assign inputArbiter_io_in_1_bits_data = feedbackOutQueue_io_deq_bits_data; // @[programmableCache.scala 242:42]
  assign inputArbiter_io_in_2_valid = io_in_otherNodes_valid; // @[programmableCache.scala 239:44]
  assign inputArbiter_io_in_2_bits_event = io_in_otherNodes_bits_event; // @[programmableCache.scala 239:44]
  assign inputArbiter_io_in_2_bits_addr = io_in_otherNodes_bits_addr; // @[programmableCache.scala 239:44]
  assign inputArbiter_io_in_2_bits_data = io_in_otherNodes_bits_data; // @[programmableCache.scala 239:44]
  assign inputArbiter_io_in_3_valid = io_in_cpu_valid; // @[programmableCache.scala 240:37]
  assign inputArbiter_io_in_3_bits_event = io_in_cpu_bits_event; // @[programmableCache.scala 240:37]
  assign inputArbiter_io_in_3_bits_addr = io_in_cpu_bits_addr; // @[programmableCache.scala 240:37]
  assign inputArbiter_io_in_3_bits_data = io_in_cpu_bits_data; // @[programmableCache.scala 240:37]
  assign inputArbiter_io_out_ready = _T_172 & _T_173; // @[programmableCache.scala 252:17]
  assign outReqArbiter_clock = clock;
  assign outReqArbiter_io_in_0_valid = reqPortQueue_0_io_deq_valid; // @[programmableCache.scala 481:41]
  assign outReqArbiter_io_in_0_bits_req_addr = reqPortQueue_0_io_deq_bits_addr; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_0_bits_req_inst = reqPortQueue_0_io_deq_bits_inst; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_0_bits_req_data = reqPortQueue_0_io_deq_bits_data; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_1_valid = reqPortQueue_1_io_deq_valid; // @[programmableCache.scala 481:41]
  assign outReqArbiter_io_in_1_bits_req_addr = reqPortQueue_1_io_deq_bits_addr; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_1_bits_req_inst = reqPortQueue_1_io_deq_bits_inst; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_1_bits_req_data = reqPortQueue_1_io_deq_bits_data; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_2_valid = reqPortQueue_2_io_deq_valid; // @[programmableCache.scala 481:41]
  assign outReqArbiter_io_in_2_bits_req_addr = reqPortQueue_2_io_deq_bits_addr; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_2_bits_req_inst = reqPortQueue_2_io_deq_bits_inst; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_2_bits_req_data = reqPortQueue_2_io_deq_bits_data; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_3_valid = reqPortQueue_3_io_deq_valid; // @[programmableCache.scala 481:41]
  assign outReqArbiter_io_in_3_bits_req_addr = reqPortQueue_3_io_deq_bits_addr; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_3_bits_req_inst = reqPortQueue_3_io_deq_bits_inst; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_3_bits_req_data = reqPortQueue_3_io_deq_bits_data; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_4_valid = reqPortQueue_4_io_deq_valid; // @[programmableCache.scala 481:41]
  assign outReqArbiter_io_in_4_bits_req_addr = reqPortQueue_4_io_deq_bits_addr; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_4_bits_req_inst = reqPortQueue_4_io_deq_bits_inst; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_4_bits_req_data = reqPortQueue_4_io_deq_bits_data; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_5_valid = reqPortQueue_5_io_deq_valid; // @[programmableCache.scala 481:41]
  assign outReqArbiter_io_in_5_bits_req_addr = reqPortQueue_5_io_deq_bits_addr; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_5_bits_req_inst = reqPortQueue_5_io_deq_bits_inst; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_5_bits_req_data = reqPortQueue_5_io_deq_bits_data; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_6_valid = reqPortQueue_6_io_deq_valid; // @[programmableCache.scala 481:41]
  assign outReqArbiter_io_in_6_bits_req_addr = reqPortQueue_6_io_deq_bits_addr; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_6_bits_req_inst = reqPortQueue_6_io_deq_bits_inst; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_6_bits_req_data = reqPortQueue_6_io_deq_bits_data; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_7_valid = reqPortQueue_7_io_deq_valid; // @[programmableCache.scala 481:41]
  assign outReqArbiter_io_in_7_bits_req_addr = reqPortQueue_7_io_deq_bits_addr; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_7_bits_req_inst = reqPortQueue_7_io_deq_bits_inst; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_7_bits_req_data = reqPortQueue_7_io_deq_bits_data; // @[programmableCache.scala 479:41]
  assign outRespArbiter_io_in_0_valid = respPortQueue_0_io_deq_valid; // @[programmableCache.scala 518:44]
  assign outRespArbiter_io_in_0_bits_addr = respPortQueue_0_io_deq_bits_addr; // @[programmableCache.scala 517:44]
  assign outRespArbiter_io_in_1_valid = respPortQueue_1_io_deq_valid; // @[programmableCache.scala 518:44]
  assign outRespArbiter_io_in_1_bits_addr = respPortQueue_1_io_deq_bits_addr; // @[programmableCache.scala 517:44]
  assign outRespArbiter_io_in_2_valid = respPortQueue_2_io_deq_valid; // @[programmableCache.scala 518:44]
  assign outRespArbiter_io_in_2_bits_addr = respPortQueue_2_io_deq_bits_addr; // @[programmableCache.scala 517:44]
  assign outRespArbiter_io_in_3_valid = respPortQueue_3_io_deq_valid; // @[programmableCache.scala 518:44]
  assign outRespArbiter_io_in_3_bits_addr = respPortQueue_3_io_deq_bits_addr; // @[programmableCache.scala 517:44]
  assign outRespArbiter_io_in_4_valid = respPortQueue_4_io_deq_valid; // @[programmableCache.scala 518:44]
  assign outRespArbiter_io_in_4_bits_addr = respPortQueue_4_io_deq_bits_addr; // @[programmableCache.scala 517:44]
  assign outRespArbiter_io_in_5_valid = respPortQueue_5_io_deq_valid; // @[programmableCache.scala 518:44]
  assign outRespArbiter_io_in_5_bits_addr = respPortQueue_5_io_deq_bits_addr; // @[programmableCache.scala 517:44]
  assign outRespArbiter_io_in_6_valid = respPortQueue_6_io_deq_valid; // @[programmableCache.scala 518:44]
  assign outRespArbiter_io_in_6_bits_addr = respPortQueue_6_io_deq_bits_addr; // @[programmableCache.scala 517:44]
  assign outRespArbiter_io_in_7_valid = respPortQueue_7_io_deq_valid; // @[programmableCache.scala 518:44]
  assign outRespArbiter_io_in_7_bits_addr = respPortQueue_7_io_deq_bits_addr; // @[programmableCache.scala 517:44]
  assign outRespArbiter_io_in_8_valid = respPortQueue_8_io_deq_valid; // @[programmableCache.scala 518:44]
  assign outRespArbiter_io_in_8_bits_addr = respPortQueue_8_io_deq_bits_addr; // @[programmableCache.scala 517:44]
  assign feedbackArbiter_io_in_0_valid = feedbackInQueue_0_io_deq_valid; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_0_bits_event = feedbackInQueue_0_io_deq_bits_event; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_0_bits_addr = feedbackInQueue_0_io_deq_bits_addr; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_0_bits_data = feedbackInQueue_0_io_deq_bits_data; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_1_valid = feedbackInQueue_1_io_deq_valid; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_1_bits_event = feedbackInQueue_1_io_deq_bits_event; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_1_bits_addr = feedbackInQueue_1_io_deq_bits_addr; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_1_bits_data = feedbackInQueue_1_io_deq_bits_data; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_2_valid = feedbackInQueue_2_io_deq_valid; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_2_bits_event = feedbackInQueue_2_io_deq_bits_event; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_2_bits_addr = feedbackInQueue_2_io_deq_bits_addr; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_2_bits_data = feedbackInQueue_2_io_deq_bits_data; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_3_valid = feedbackInQueue_3_io_deq_valid; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_3_bits_event = feedbackInQueue_3_io_deq_bits_event; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_3_bits_addr = feedbackInQueue_3_io_deq_bits_addr; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_3_bits_data = feedbackInQueue_3_io_deq_bits_data; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_4_valid = feedbackInQueue_4_io_deq_valid; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_4_bits_event = feedbackInQueue_4_io_deq_bits_event; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_4_bits_addr = feedbackInQueue_4_io_deq_bits_addr; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_4_bits_data = feedbackInQueue_4_io_deq_bits_data; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_5_valid = feedbackInQueue_5_io_deq_valid; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_5_bits_event = feedbackInQueue_5_io_deq_bits_event; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_5_bits_addr = feedbackInQueue_5_io_deq_bits_addr; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_5_bits_data = feedbackInQueue_5_io_deq_bits_data; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_6_valid = feedbackInQueue_6_io_deq_valid; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_6_bits_event = feedbackInQueue_6_io_deq_bits_event; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_6_bits_addr = feedbackInQueue_6_io_deq_bits_addr; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_6_bits_data = feedbackInQueue_6_io_deq_bits_data; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_7_valid = feedbackInQueue_7_io_deq_valid; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_7_bits_event = feedbackInQueue_7_io_deq_bits_event; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_7_bits_addr = feedbackInQueue_7_io_deq_bits_addr; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_7_bits_data = feedbackInQueue_7_io_deq_bits_data; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_out_ready = feedbackOutQueue_io_enq_ready; // @[programmableCache.scala 244:29]
  assign input__clock = clock;
  assign input__reset = reset;
  assign input__io_enq_valid = _T_178 & _T_173; // @[programmableCache.scala 286:24]
  assign input__io_enq_bits_inst_event = inputArbiter_io_out_bits_event; // @[programmableCache.scala 288:28]
  assign input__io_enq_bits_inst_addr = inputArbiter_io_out_bits_addr; // @[programmableCache.scala 288:28]
  assign input__io_enq_bits_inst_data = inputArbiter_io_out_bits_data; // @[programmableCache.scala 288:28]
  assign input__io_enq_bits_tbeOut_state_state = tbe_io_outputTBE_bits_state_state; // @[programmableCache.scala 289:30]
  assign input__io_enq_bits_tbeOut_way = tbe_io_outputTBE_bits_way; // @[programmableCache.scala 289:30]
  assign input__io_enq_bits_tbeOut_fields_0 = tbe_io_outputTBE_bits_fields_0; // @[programmableCache.scala 289:30]
  assign input__io_deq_ready = routineQueue_io_enq_ready; // @[programmableCache.scala 351:24]
  assign respPortQueue_0_clock = clock;
  assign respPortQueue_0_reset = reset;
  assign respPortQueue_0_io_enq_valid = cache_io_cpu_0_resp_valid & cache_io_cpu_0_resp_bits_iswrite; // @[programmableCache.scala 506:44]
  assign respPortQueue_0_io_enq_bits_event = 2'h0; // @[programmableCache.scala 504:44]
  assign respPortQueue_0_io_enq_bits_addr = actionReg_0_io_deq_bits_addr; // @[programmableCache.scala 505:44]
  assign respPortQueue_0_io_enq_bits_data = 64'h0; // @[programmableCache.scala 503:44]
  assign respPortQueue_0_io_deq_ready = 1'h1; // @[programmableCache.scala 519:39]
  assign respPortQueue_1_clock = clock;
  assign respPortQueue_1_reset = reset;
  assign respPortQueue_1_io_enq_valid = cache_io_cpu_1_resp_valid & cache_io_cpu_1_resp_bits_iswrite; // @[programmableCache.scala 506:44]
  assign respPortQueue_1_io_enq_bits_event = 2'h0; // @[programmableCache.scala 504:44]
  assign respPortQueue_1_io_enq_bits_addr = actionReg_1_io_deq_bits_addr; // @[programmableCache.scala 505:44]
  assign respPortQueue_1_io_enq_bits_data = 64'h0; // @[programmableCache.scala 503:44]
  assign respPortQueue_1_io_deq_ready = 1'h1; // @[programmableCache.scala 519:39]
  assign respPortQueue_2_clock = clock;
  assign respPortQueue_2_reset = reset;
  assign respPortQueue_2_io_enq_valid = cache_io_cpu_2_resp_valid & cache_io_cpu_2_resp_bits_iswrite; // @[programmableCache.scala 506:44]
  assign respPortQueue_2_io_enq_bits_event = 2'h0; // @[programmableCache.scala 504:44]
  assign respPortQueue_2_io_enq_bits_addr = actionReg_2_io_deq_bits_addr; // @[programmableCache.scala 505:44]
  assign respPortQueue_2_io_enq_bits_data = 64'h0; // @[programmableCache.scala 503:44]
  assign respPortQueue_2_io_deq_ready = 1'h1; // @[programmableCache.scala 519:39]
  assign respPortQueue_3_clock = clock;
  assign respPortQueue_3_reset = reset;
  assign respPortQueue_3_io_enq_valid = cache_io_cpu_3_resp_valid & cache_io_cpu_3_resp_bits_iswrite; // @[programmableCache.scala 506:44]
  assign respPortQueue_3_io_enq_bits_event = 2'h0; // @[programmableCache.scala 504:44]
  assign respPortQueue_3_io_enq_bits_addr = actionReg_3_io_deq_bits_addr; // @[programmableCache.scala 505:44]
  assign respPortQueue_3_io_enq_bits_data = 64'h0; // @[programmableCache.scala 503:44]
  assign respPortQueue_3_io_deq_ready = 1'h1; // @[programmableCache.scala 519:39]
  assign respPortQueue_4_clock = clock;
  assign respPortQueue_4_reset = reset;
  assign respPortQueue_4_io_enq_valid = cache_io_cpu_4_resp_valid & cache_io_cpu_4_resp_bits_iswrite; // @[programmableCache.scala 506:44]
  assign respPortQueue_4_io_enq_bits_event = 2'h0; // @[programmableCache.scala 504:44]
  assign respPortQueue_4_io_enq_bits_addr = actionReg_4_io_deq_bits_addr; // @[programmableCache.scala 505:44]
  assign respPortQueue_4_io_enq_bits_data = 64'h0; // @[programmableCache.scala 503:44]
  assign respPortQueue_4_io_deq_ready = 1'h1; // @[programmableCache.scala 519:39]
  assign respPortQueue_5_clock = clock;
  assign respPortQueue_5_reset = reset;
  assign respPortQueue_5_io_enq_valid = cache_io_cpu_5_resp_valid & cache_io_cpu_5_resp_bits_iswrite; // @[programmableCache.scala 506:44]
  assign respPortQueue_5_io_enq_bits_event = 2'h0; // @[programmableCache.scala 504:44]
  assign respPortQueue_5_io_enq_bits_addr = actionReg_5_io_deq_bits_addr; // @[programmableCache.scala 505:44]
  assign respPortQueue_5_io_enq_bits_data = 64'h0; // @[programmableCache.scala 503:44]
  assign respPortQueue_5_io_deq_ready = 1'h1; // @[programmableCache.scala 519:39]
  assign respPortQueue_6_clock = clock;
  assign respPortQueue_6_reset = reset;
  assign respPortQueue_6_io_enq_valid = cache_io_cpu_6_resp_valid & cache_io_cpu_6_resp_bits_iswrite; // @[programmableCache.scala 506:44]
  assign respPortQueue_6_io_enq_bits_event = 2'h0; // @[programmableCache.scala 504:44]
  assign respPortQueue_6_io_enq_bits_addr = actionReg_6_io_deq_bits_addr; // @[programmableCache.scala 505:44]
  assign respPortQueue_6_io_enq_bits_data = 64'h0; // @[programmableCache.scala 503:44]
  assign respPortQueue_6_io_deq_ready = 1'h1; // @[programmableCache.scala 519:39]
  assign respPortQueue_7_clock = clock;
  assign respPortQueue_7_reset = reset;
  assign respPortQueue_7_io_enq_valid = cache_io_cpu_7_resp_valid & cache_io_cpu_7_resp_bits_iswrite; // @[programmableCache.scala 506:44]
  assign respPortQueue_7_io_enq_bits_event = 2'h0; // @[programmableCache.scala 504:44]
  assign respPortQueue_7_io_enq_bits_addr = actionReg_7_io_deq_bits_addr; // @[programmableCache.scala 505:44]
  assign respPortQueue_7_io_enq_bits_data = 64'h0; // @[programmableCache.scala 503:44]
  assign respPortQueue_7_io_deq_ready = 1'h1; // @[programmableCache.scala 519:39]
  assign respPortQueue_8_clock = clock;
  assign respPortQueue_8_reset = reset;
  assign respPortQueue_8_io_enq_valid = cache_io_bipassLD_out_valid; // @[programmableCache.scala 512:45]
  assign respPortQueue_8_io_enq_bits_event = 2'h0; // @[programmableCache.scala 510:45]
  assign respPortQueue_8_io_enq_bits_addr = _T_783; // @[programmableCache.scala 511:45]
  assign respPortQueue_8_io_enq_bits_data = cache_io_bipassLD_out_bits_data; // @[programmableCache.scala 509:45]
  assign respPortQueue_8_io_deq_ready = 1'h1; // @[programmableCache.scala 519:39]
  assign reqPortQueue_0_clock = clock;
  assign reqPortQueue_0_reset = reset;
  assign reqPortQueue_0_io_enq_valid = _T_282 & actionReg_0_io_deq_valid; // @[programmableCache.scala 490:38]
  assign reqPortQueue_0_io_enq_bits_addr = actionReg_0_io_deq_bits_addr; // @[programmableCache.scala 488:42]
  assign reqPortQueue_0_io_enq_bits_inst = 8'h0; // @[programmableCache.scala 489:41]
  assign reqPortQueue_0_io_enq_bits_data = actionReg_0_io_deq_bits_action_signals[0] ? _GEN_1481 : {{32'd0}, actionReg_0_io_deq_bits_addr}; // @[programmableCache.scala 487:41]
  assign reqPortQueue_0_io_deq_ready = outReqArbiter_io_in_0_ready; // @[programmableCache.scala 482:38]
  assign reqPortQueue_1_clock = clock;
  assign reqPortQueue_1_reset = reset;
  assign reqPortQueue_1_io_enq_valid = _T_339 & actionReg_1_io_deq_valid; // @[programmableCache.scala 490:38]
  assign reqPortQueue_1_io_enq_bits_addr = actionReg_1_io_deq_bits_addr; // @[programmableCache.scala 488:42]
  assign reqPortQueue_1_io_enq_bits_inst = 8'h0; // @[programmableCache.scala 489:41]
  assign reqPortQueue_1_io_enq_bits_data = actionReg_1_io_deq_bits_action_signals[0] ? _GEN_1485 : {{32'd0}, actionReg_1_io_deq_bits_addr}; // @[programmableCache.scala 487:41]
  assign reqPortQueue_1_io_deq_ready = outReqArbiter_io_in_1_ready; // @[programmableCache.scala 482:38]
  assign reqPortQueue_2_clock = clock;
  assign reqPortQueue_2_reset = reset;
  assign reqPortQueue_2_io_enq_valid = _T_396 & actionReg_2_io_deq_valid; // @[programmableCache.scala 490:38]
  assign reqPortQueue_2_io_enq_bits_addr = actionReg_2_io_deq_bits_addr; // @[programmableCache.scala 488:42]
  assign reqPortQueue_2_io_enq_bits_inst = 8'h0; // @[programmableCache.scala 489:41]
  assign reqPortQueue_2_io_enq_bits_data = actionReg_2_io_deq_bits_action_signals[0] ? _GEN_1489 : {{32'd0}, actionReg_2_io_deq_bits_addr}; // @[programmableCache.scala 487:41]
  assign reqPortQueue_2_io_deq_ready = outReqArbiter_io_in_2_ready; // @[programmableCache.scala 482:38]
  assign reqPortQueue_3_clock = clock;
  assign reqPortQueue_3_reset = reset;
  assign reqPortQueue_3_io_enq_valid = _T_453 & actionReg_3_io_deq_valid; // @[programmableCache.scala 490:38]
  assign reqPortQueue_3_io_enq_bits_addr = actionReg_3_io_deq_bits_addr; // @[programmableCache.scala 488:42]
  assign reqPortQueue_3_io_enq_bits_inst = 8'h0; // @[programmableCache.scala 489:41]
  assign reqPortQueue_3_io_enq_bits_data = actionReg_3_io_deq_bits_action_signals[0] ? _GEN_1493 : {{32'd0}, actionReg_3_io_deq_bits_addr}; // @[programmableCache.scala 487:41]
  assign reqPortQueue_3_io_deq_ready = outReqArbiter_io_in_3_ready; // @[programmableCache.scala 482:38]
  assign reqPortQueue_4_clock = clock;
  assign reqPortQueue_4_reset = reset;
  assign reqPortQueue_4_io_enq_valid = _T_510 & actionReg_4_io_deq_valid; // @[programmableCache.scala 490:38]
  assign reqPortQueue_4_io_enq_bits_addr = actionReg_4_io_deq_bits_addr; // @[programmableCache.scala 488:42]
  assign reqPortQueue_4_io_enq_bits_inst = 8'h0; // @[programmableCache.scala 489:41]
  assign reqPortQueue_4_io_enq_bits_data = actionReg_4_io_deq_bits_action_signals[0] ? _GEN_1497 : {{32'd0}, actionReg_4_io_deq_bits_addr}; // @[programmableCache.scala 487:41]
  assign reqPortQueue_4_io_deq_ready = outReqArbiter_io_in_4_ready; // @[programmableCache.scala 482:38]
  assign reqPortQueue_5_clock = clock;
  assign reqPortQueue_5_reset = reset;
  assign reqPortQueue_5_io_enq_valid = _T_567 & actionReg_5_io_deq_valid; // @[programmableCache.scala 490:38]
  assign reqPortQueue_5_io_enq_bits_addr = actionReg_5_io_deq_bits_addr; // @[programmableCache.scala 488:42]
  assign reqPortQueue_5_io_enq_bits_inst = 8'h0; // @[programmableCache.scala 489:41]
  assign reqPortQueue_5_io_enq_bits_data = actionReg_5_io_deq_bits_action_signals[0] ? _GEN_1501 : {{32'd0}, actionReg_5_io_deq_bits_addr}; // @[programmableCache.scala 487:41]
  assign reqPortQueue_5_io_deq_ready = outReqArbiter_io_in_5_ready; // @[programmableCache.scala 482:38]
  assign reqPortQueue_6_clock = clock;
  assign reqPortQueue_6_reset = reset;
  assign reqPortQueue_6_io_enq_valid = _T_624 & actionReg_6_io_deq_valid; // @[programmableCache.scala 490:38]
  assign reqPortQueue_6_io_enq_bits_addr = actionReg_6_io_deq_bits_addr; // @[programmableCache.scala 488:42]
  assign reqPortQueue_6_io_enq_bits_inst = 8'h0; // @[programmableCache.scala 489:41]
  assign reqPortQueue_6_io_enq_bits_data = actionReg_6_io_deq_bits_action_signals[0] ? _GEN_1505 : {{32'd0}, actionReg_6_io_deq_bits_addr}; // @[programmableCache.scala 487:41]
  assign reqPortQueue_6_io_deq_ready = outReqArbiter_io_in_6_ready; // @[programmableCache.scala 482:38]
  assign reqPortQueue_7_clock = clock;
  assign reqPortQueue_7_reset = reset;
  assign reqPortQueue_7_io_enq_valid = _T_681 & actionReg_7_io_deq_valid; // @[programmableCache.scala 490:38]
  assign reqPortQueue_7_io_enq_bits_addr = actionReg_7_io_deq_bits_addr; // @[programmableCache.scala 488:42]
  assign reqPortQueue_7_io_enq_bits_inst = 8'h0; // @[programmableCache.scala 489:41]
  assign reqPortQueue_7_io_enq_bits_data = actionReg_7_io_deq_bits_action_signals[0] ? _GEN_1509 : {{32'd0}, actionReg_7_io_deq_bits_addr}; // @[programmableCache.scala 487:41]
  assign reqPortQueue_7_io_deq_ready = outReqArbiter_io_in_7_ready; // @[programmableCache.scala 482:38]
  assign feedbackInQueue_0_clock = clock;
  assign feedbackInQueue_0_reset = reset;
  assign feedbackInQueue_0_io_enq_valid = _T_278 & actionReg_0_io_deq_valid; // @[programmableCache.scala 250:41]
  assign feedbackInQueue_0_io_enq_bits_event = actionReg_0_io_deq_bits_action_signals[13:12]; // @[programmableCache.scala 248:46]
  assign feedbackInQueue_0_io_enq_bits_addr = actionReg_0_io_deq_bits_addr + _GEN_1510; // @[programmableCache.scala 247:45]
  assign feedbackInQueue_0_io_enq_bits_data = actionReg_0_io_deq_bits_data - _GEN_1511; // @[programmableCache.scala 249:45]
  assign feedbackInQueue_0_io_deq_ready = feedbackArbiter_io_in_0_ready; // @[programmableCache.scala 246:34]
  assign feedbackInQueue_1_clock = clock;
  assign feedbackInQueue_1_reset = reset;
  assign feedbackInQueue_1_io_enq_valid = _T_335 & actionReg_1_io_deq_valid; // @[programmableCache.scala 250:41]
  assign feedbackInQueue_1_io_enq_bits_event = actionReg_1_io_deq_bits_action_signals[13:12]; // @[programmableCache.scala 248:46]
  assign feedbackInQueue_1_io_enq_bits_addr = actionReg_1_io_deq_bits_addr + _GEN_1512; // @[programmableCache.scala 247:45]
  assign feedbackInQueue_1_io_enq_bits_data = actionReg_1_io_deq_bits_data - _GEN_1513; // @[programmableCache.scala 249:45]
  assign feedbackInQueue_1_io_deq_ready = feedbackArbiter_io_in_1_ready; // @[programmableCache.scala 246:34]
  assign feedbackInQueue_2_clock = clock;
  assign feedbackInQueue_2_reset = reset;
  assign feedbackInQueue_2_io_enq_valid = _T_392 & actionReg_2_io_deq_valid; // @[programmableCache.scala 250:41]
  assign feedbackInQueue_2_io_enq_bits_event = actionReg_2_io_deq_bits_action_signals[13:12]; // @[programmableCache.scala 248:46]
  assign feedbackInQueue_2_io_enq_bits_addr = actionReg_2_io_deq_bits_addr + _GEN_1514; // @[programmableCache.scala 247:45]
  assign feedbackInQueue_2_io_enq_bits_data = actionReg_2_io_deq_bits_data - _GEN_1515; // @[programmableCache.scala 249:45]
  assign feedbackInQueue_2_io_deq_ready = feedbackArbiter_io_in_2_ready; // @[programmableCache.scala 246:34]
  assign feedbackInQueue_3_clock = clock;
  assign feedbackInQueue_3_reset = reset;
  assign feedbackInQueue_3_io_enq_valid = _T_449 & actionReg_3_io_deq_valid; // @[programmableCache.scala 250:41]
  assign feedbackInQueue_3_io_enq_bits_event = actionReg_3_io_deq_bits_action_signals[13:12]; // @[programmableCache.scala 248:46]
  assign feedbackInQueue_3_io_enq_bits_addr = actionReg_3_io_deq_bits_addr + _GEN_1516; // @[programmableCache.scala 247:45]
  assign feedbackInQueue_3_io_enq_bits_data = actionReg_3_io_deq_bits_data - _GEN_1517; // @[programmableCache.scala 249:45]
  assign feedbackInQueue_3_io_deq_ready = feedbackArbiter_io_in_3_ready; // @[programmableCache.scala 246:34]
  assign feedbackInQueue_4_clock = clock;
  assign feedbackInQueue_4_reset = reset;
  assign feedbackInQueue_4_io_enq_valid = _T_506 & actionReg_4_io_deq_valid; // @[programmableCache.scala 250:41]
  assign feedbackInQueue_4_io_enq_bits_event = actionReg_4_io_deq_bits_action_signals[13:12]; // @[programmableCache.scala 248:46]
  assign feedbackInQueue_4_io_enq_bits_addr = actionReg_4_io_deq_bits_addr + _GEN_1518; // @[programmableCache.scala 247:45]
  assign feedbackInQueue_4_io_enq_bits_data = actionReg_4_io_deq_bits_data - _GEN_1519; // @[programmableCache.scala 249:45]
  assign feedbackInQueue_4_io_deq_ready = feedbackArbiter_io_in_4_ready; // @[programmableCache.scala 246:34]
  assign feedbackInQueue_5_clock = clock;
  assign feedbackInQueue_5_reset = reset;
  assign feedbackInQueue_5_io_enq_valid = _T_563 & actionReg_5_io_deq_valid; // @[programmableCache.scala 250:41]
  assign feedbackInQueue_5_io_enq_bits_event = actionReg_5_io_deq_bits_action_signals[13:12]; // @[programmableCache.scala 248:46]
  assign feedbackInQueue_5_io_enq_bits_addr = actionReg_5_io_deq_bits_addr + _GEN_1520; // @[programmableCache.scala 247:45]
  assign feedbackInQueue_5_io_enq_bits_data = actionReg_5_io_deq_bits_data - _GEN_1521; // @[programmableCache.scala 249:45]
  assign feedbackInQueue_5_io_deq_ready = feedbackArbiter_io_in_5_ready; // @[programmableCache.scala 246:34]
  assign feedbackInQueue_6_clock = clock;
  assign feedbackInQueue_6_reset = reset;
  assign feedbackInQueue_6_io_enq_valid = _T_620 & actionReg_6_io_deq_valid; // @[programmableCache.scala 250:41]
  assign feedbackInQueue_6_io_enq_bits_event = actionReg_6_io_deq_bits_action_signals[13:12]; // @[programmableCache.scala 248:46]
  assign feedbackInQueue_6_io_enq_bits_addr = actionReg_6_io_deq_bits_addr + _GEN_1522; // @[programmableCache.scala 247:45]
  assign feedbackInQueue_6_io_enq_bits_data = actionReg_6_io_deq_bits_data - _GEN_1523; // @[programmableCache.scala 249:45]
  assign feedbackInQueue_6_io_deq_ready = feedbackArbiter_io_in_6_ready; // @[programmableCache.scala 246:34]
  assign feedbackInQueue_7_clock = clock;
  assign feedbackInQueue_7_reset = reset;
  assign feedbackInQueue_7_io_enq_valid = _T_677 & actionReg_7_io_deq_valid; // @[programmableCache.scala 250:41]
  assign feedbackInQueue_7_io_enq_bits_event = actionReg_7_io_deq_bits_action_signals[13:12]; // @[programmableCache.scala 248:46]
  assign feedbackInQueue_7_io_enq_bits_addr = actionReg_7_io_deq_bits_addr + _GEN_1524; // @[programmableCache.scala 247:45]
  assign feedbackInQueue_7_io_enq_bits_data = actionReg_7_io_deq_bits_data - _GEN_1525; // @[programmableCache.scala 249:45]
  assign feedbackInQueue_7_io_deq_ready = feedbackArbiter_io_in_7_ready; // @[programmableCache.scala 246:34]
  assign probeWay_clock = clock;
  assign probeWay_reset = reset;
  assign probeWay_io_enq_valid = cache_io_probe_resp_valid; // @[programmableCache.scala 217:29]
  assign probeWay_io_enq_bits = cache_io_probe_resp_bits_way; // @[programmableCache.scala 216:28]
  assign probeWay_io_deq_ready = input__io_deq_ready & input__io_deq_valid; // @[programmableCache.scala 227:29]
  assign feedbackOutQueue_clock = clock;
  assign feedbackOutQueue_reset = reset;
  assign feedbackOutQueue_io_enq_valid = feedbackArbiter_io_out_valid; // @[programmableCache.scala 244:29]
  assign feedbackOutQueue_io_enq_bits_event = feedbackArbiter_io_out_bits_event; // @[programmableCache.scala 244:29]
  assign feedbackOutQueue_io_enq_bits_addr = feedbackArbiter_io_out_bits_addr; // @[programmableCache.scala 244:29]
  assign feedbackOutQueue_io_enq_bits_data = feedbackArbiter_io_out_bits_data; // @[programmableCache.scala 244:29]
  assign feedbackOutQueue_io_deq_ready = inputArbiter_io_in_1_ready; // @[programmableCache.scala 242:42]
  assign routineQueue_clock = clock;
  assign routineQueue_reset = reset;
  assign routineQueue_io_enq_valid = input__io_deq_valid; // @[programmableCache.scala 350:31]
  assign routineQueue_io_enq_bits = {{10'd0}, _GEN_15}; // @[programmableCache.scala 349:30]
  assign routineQueue_io_deq_ready = ~pc_io_isFull; // @[programmableCache.scala 352:31]
  assign actionReg_0_clock = clock;
  assign actionReg_0_reset = reset;
  assign actionReg_0_io_enq_valid = pc_io_read_0_out_bits_valid; // @[programmableCache.scala 438:35]
  assign actionReg_0_io_enq_bits_addr = pc_io_read_0_out_bits_addr; // @[programmableCache.scala 385:39]
  assign actionReg_0_io_enq_bits_way = _T_290[1:0]; // @[programmableCache.scala 386:39]
  assign actionReg_0_io_enq_bits_data = pc_io_read_0_out_bits_data; // @[programmableCache.scala 387:39]
  assign actionReg_0_io_enq_bits_replaceWay = pc_io_read_0_out_bits_replaceWay; // @[programmableCache.scala 388:45]
  assign actionReg_0_io_enq_bits_tbeFields_0 = pc_io_read_0_out_bits_tbeFields_0; // @[programmableCache.scala 390:44]
  assign actionReg_0_io_enq_bits_action_signals = _GEN_88[27:0]; // @[programmableCache.scala 383:49]
  assign actionReg_0_io_enq_bits_action_actionType = _GEN_88[31:28]; // @[programmableCache.scala 384:52]
  assign actionReg_0_io_deq_ready = 1'h1; // @[programmableCache.scala 437:35]
  assign actionReg_1_clock = clock;
  assign actionReg_1_reset = reset;
  assign actionReg_1_io_enq_valid = pc_io_read_1_out_bits_valid; // @[programmableCache.scala 438:35]
  assign actionReg_1_io_enq_bits_addr = pc_io_read_1_out_bits_addr; // @[programmableCache.scala 385:39]
  assign actionReg_1_io_enq_bits_way = _T_347[1:0]; // @[programmableCache.scala 386:39]
  assign actionReg_1_io_enq_bits_data = pc_io_read_1_out_bits_data; // @[programmableCache.scala 387:39]
  assign actionReg_1_io_enq_bits_replaceWay = pc_io_read_1_out_bits_replaceWay; // @[programmableCache.scala 388:45]
  assign actionReg_1_io_enq_bits_tbeFields_0 = pc_io_read_1_out_bits_tbeFields_0; // @[programmableCache.scala 390:44]
  assign actionReg_1_io_enq_bits_action_signals = _GEN_269[27:0]; // @[programmableCache.scala 383:49]
  assign actionReg_1_io_enq_bits_action_actionType = _GEN_269[31:28]; // @[programmableCache.scala 384:52]
  assign actionReg_1_io_deq_ready = 1'h1; // @[programmableCache.scala 437:35]
  assign actionReg_2_clock = clock;
  assign actionReg_2_reset = reset;
  assign actionReg_2_io_enq_valid = pc_io_read_2_out_bits_valid; // @[programmableCache.scala 438:35]
  assign actionReg_2_io_enq_bits_addr = pc_io_read_2_out_bits_addr; // @[programmableCache.scala 385:39]
  assign actionReg_2_io_enq_bits_way = _T_404[1:0]; // @[programmableCache.scala 386:39]
  assign actionReg_2_io_enq_bits_data = pc_io_read_2_out_bits_data; // @[programmableCache.scala 387:39]
  assign actionReg_2_io_enq_bits_replaceWay = pc_io_read_2_out_bits_replaceWay; // @[programmableCache.scala 388:45]
  assign actionReg_2_io_enq_bits_tbeFields_0 = pc_io_read_2_out_bits_tbeFields_0; // @[programmableCache.scala 390:44]
  assign actionReg_2_io_enq_bits_action_signals = _GEN_450[27:0]; // @[programmableCache.scala 383:49]
  assign actionReg_2_io_enq_bits_action_actionType = _GEN_450[31:28]; // @[programmableCache.scala 384:52]
  assign actionReg_2_io_deq_ready = 1'h1; // @[programmableCache.scala 437:35]
  assign actionReg_3_clock = clock;
  assign actionReg_3_reset = reset;
  assign actionReg_3_io_enq_valid = pc_io_read_3_out_bits_valid; // @[programmableCache.scala 438:35]
  assign actionReg_3_io_enq_bits_addr = pc_io_read_3_out_bits_addr; // @[programmableCache.scala 385:39]
  assign actionReg_3_io_enq_bits_way = _T_461[1:0]; // @[programmableCache.scala 386:39]
  assign actionReg_3_io_enq_bits_data = pc_io_read_3_out_bits_data; // @[programmableCache.scala 387:39]
  assign actionReg_3_io_enq_bits_replaceWay = pc_io_read_3_out_bits_replaceWay; // @[programmableCache.scala 388:45]
  assign actionReg_3_io_enq_bits_tbeFields_0 = pc_io_read_3_out_bits_tbeFields_0; // @[programmableCache.scala 390:44]
  assign actionReg_3_io_enq_bits_action_signals = _GEN_631[27:0]; // @[programmableCache.scala 383:49]
  assign actionReg_3_io_enq_bits_action_actionType = _GEN_631[31:28]; // @[programmableCache.scala 384:52]
  assign actionReg_3_io_deq_ready = 1'h1; // @[programmableCache.scala 437:35]
  assign actionReg_4_clock = clock;
  assign actionReg_4_reset = reset;
  assign actionReg_4_io_enq_valid = pc_io_read_4_out_bits_valid; // @[programmableCache.scala 438:35]
  assign actionReg_4_io_enq_bits_addr = pc_io_read_4_out_bits_addr; // @[programmableCache.scala 385:39]
  assign actionReg_4_io_enq_bits_way = _T_518[1:0]; // @[programmableCache.scala 386:39]
  assign actionReg_4_io_enq_bits_data = pc_io_read_4_out_bits_data; // @[programmableCache.scala 387:39]
  assign actionReg_4_io_enq_bits_replaceWay = pc_io_read_4_out_bits_replaceWay; // @[programmableCache.scala 388:45]
  assign actionReg_4_io_enq_bits_tbeFields_0 = pc_io_read_4_out_bits_tbeFields_0; // @[programmableCache.scala 390:44]
  assign actionReg_4_io_enq_bits_action_signals = _GEN_812[27:0]; // @[programmableCache.scala 383:49]
  assign actionReg_4_io_enq_bits_action_actionType = _GEN_812[31:28]; // @[programmableCache.scala 384:52]
  assign actionReg_4_io_deq_ready = 1'h1; // @[programmableCache.scala 437:35]
  assign actionReg_5_clock = clock;
  assign actionReg_5_reset = reset;
  assign actionReg_5_io_enq_valid = pc_io_read_5_out_bits_valid; // @[programmableCache.scala 438:35]
  assign actionReg_5_io_enq_bits_addr = pc_io_read_5_out_bits_addr; // @[programmableCache.scala 385:39]
  assign actionReg_5_io_enq_bits_way = _T_575[1:0]; // @[programmableCache.scala 386:39]
  assign actionReg_5_io_enq_bits_data = pc_io_read_5_out_bits_data; // @[programmableCache.scala 387:39]
  assign actionReg_5_io_enq_bits_replaceWay = pc_io_read_5_out_bits_replaceWay; // @[programmableCache.scala 388:45]
  assign actionReg_5_io_enq_bits_tbeFields_0 = pc_io_read_5_out_bits_tbeFields_0; // @[programmableCache.scala 390:44]
  assign actionReg_5_io_enq_bits_action_signals = _GEN_993[27:0]; // @[programmableCache.scala 383:49]
  assign actionReg_5_io_enq_bits_action_actionType = _GEN_993[31:28]; // @[programmableCache.scala 384:52]
  assign actionReg_5_io_deq_ready = 1'h1; // @[programmableCache.scala 437:35]
  assign actionReg_6_clock = clock;
  assign actionReg_6_reset = reset;
  assign actionReg_6_io_enq_valid = pc_io_read_6_out_bits_valid; // @[programmableCache.scala 438:35]
  assign actionReg_6_io_enq_bits_addr = pc_io_read_6_out_bits_addr; // @[programmableCache.scala 385:39]
  assign actionReg_6_io_enq_bits_way = _T_632[1:0]; // @[programmableCache.scala 386:39]
  assign actionReg_6_io_enq_bits_data = pc_io_read_6_out_bits_data; // @[programmableCache.scala 387:39]
  assign actionReg_6_io_enq_bits_replaceWay = pc_io_read_6_out_bits_replaceWay; // @[programmableCache.scala 388:45]
  assign actionReg_6_io_enq_bits_tbeFields_0 = pc_io_read_6_out_bits_tbeFields_0; // @[programmableCache.scala 390:44]
  assign actionReg_6_io_enq_bits_action_signals = _GEN_1174[27:0]; // @[programmableCache.scala 383:49]
  assign actionReg_6_io_enq_bits_action_actionType = _GEN_1174[31:28]; // @[programmableCache.scala 384:52]
  assign actionReg_6_io_deq_ready = 1'h1; // @[programmableCache.scala 437:35]
  assign actionReg_7_clock = clock;
  assign actionReg_7_reset = reset;
  assign actionReg_7_io_enq_valid = pc_io_read_7_out_bits_valid; // @[programmableCache.scala 438:35]
  assign actionReg_7_io_enq_bits_addr = pc_io_read_7_out_bits_addr; // @[programmableCache.scala 385:39]
  assign actionReg_7_io_enq_bits_way = _T_689[1:0]; // @[programmableCache.scala 386:39]
  assign actionReg_7_io_enq_bits_data = pc_io_read_7_out_bits_data; // @[programmableCache.scala 387:39]
  assign actionReg_7_io_enq_bits_replaceWay = pc_io_read_7_out_bits_replaceWay; // @[programmableCache.scala 388:45]
  assign actionReg_7_io_enq_bits_tbeFields_0 = pc_io_read_7_out_bits_tbeFields_0; // @[programmableCache.scala 390:44]
  assign actionReg_7_io_enq_bits_action_signals = _GEN_1355[27:0]; // @[programmableCache.scala 383:49]
  assign actionReg_7_io_enq_bits_action_actionType = _GEN_1355[31:28]; // @[programmableCache.scala 384:52]
  assign actionReg_7_io_deq_ready = 1'h1; // @[programmableCache.scala 437:35]
  assign mimoQ_clock = clock;
  assign mimoQ_reset = reset;
  assign mimoQ_io_enq_valid = cache_io_probe_multiWay_valid; // @[programmableCache.scala 222:24]
  assign mimoQ_io_enq_bits_0_way = cache_io_probe_multiWay_bits_way_0; // @[programmableCache.scala 219:56]
  assign mimoQ_io_enq_bits_0_addr = cache_io_probe_multiWay_bits_addr; // @[programmableCache.scala 220:57]
  assign mimoQ_io_enq_bits_1_way = cache_io_probe_multiWay_bits_way_1; // @[programmableCache.scala 219:56]
  assign mimoQ_io_enq_bits_1_addr = cache_io_probe_multiWay_bits_addr; // @[programmableCache.scala 220:57]
  assign compUnit_0_clock = clock;
  assign compUnit_0_reset = reset;
  assign compUnit_0_io_instruction_valid = _T_284 & actionReg_0_io_deq_valid; // @[programmableCache.scala 435:42]
  assign compUnit_0_io_instruction_bits = actionReg_0_io_deq_bits_action_signals; // @[programmableCache.scala 434:41]
  assign compUnit_0_io_clear = _T_280 & actionReg_0_io_deq_valid; // @[programmableCache.scala 381:30]
  assign compUnit_0_io_op1_valid = compUnitInput1_0_io_out_valid; // @[programmableCache.scala 425:28]
  assign compUnit_0_io_op1_bits = compUnitInput1_0_io_out_bits; // @[programmableCache.scala 425:28]
  assign compUnit_0_io_op2_valid = compUnitInput2_0_io_out_valid; // @[programmableCache.scala 432:28]
  assign compUnit_0_io_op2_bits = compUnitInput2_0_io_out_bits; // @[programmableCache.scala 432:28]
  assign compUnit_1_clock = clock;
  assign compUnit_1_reset = reset;
  assign compUnit_1_io_instruction_valid = _T_341 & actionReg_1_io_deq_valid; // @[programmableCache.scala 435:42]
  assign compUnit_1_io_instruction_bits = actionReg_1_io_deq_bits_action_signals; // @[programmableCache.scala 434:41]
  assign compUnit_1_io_clear = _T_337 & actionReg_1_io_deq_valid; // @[programmableCache.scala 381:30]
  assign compUnit_1_io_op1_valid = compUnitInput1_1_io_out_valid; // @[programmableCache.scala 425:28]
  assign compUnit_1_io_op1_bits = compUnitInput1_1_io_out_bits; // @[programmableCache.scala 425:28]
  assign compUnit_1_io_op2_valid = compUnitInput2_1_io_out_valid; // @[programmableCache.scala 432:28]
  assign compUnit_1_io_op2_bits = compUnitInput2_1_io_out_bits; // @[programmableCache.scala 432:28]
  assign compUnit_2_clock = clock;
  assign compUnit_2_reset = reset;
  assign compUnit_2_io_instruction_valid = _T_398 & actionReg_2_io_deq_valid; // @[programmableCache.scala 435:42]
  assign compUnit_2_io_instruction_bits = actionReg_2_io_deq_bits_action_signals; // @[programmableCache.scala 434:41]
  assign compUnit_2_io_clear = _T_394 & actionReg_2_io_deq_valid; // @[programmableCache.scala 381:30]
  assign compUnit_2_io_op1_valid = compUnitInput1_2_io_out_valid; // @[programmableCache.scala 425:28]
  assign compUnit_2_io_op1_bits = compUnitInput1_2_io_out_bits; // @[programmableCache.scala 425:28]
  assign compUnit_2_io_op2_valid = compUnitInput2_2_io_out_valid; // @[programmableCache.scala 432:28]
  assign compUnit_2_io_op2_bits = compUnitInput2_2_io_out_bits; // @[programmableCache.scala 432:28]
  assign compUnit_3_clock = clock;
  assign compUnit_3_reset = reset;
  assign compUnit_3_io_instruction_valid = _T_455 & actionReg_3_io_deq_valid; // @[programmableCache.scala 435:42]
  assign compUnit_3_io_instruction_bits = actionReg_3_io_deq_bits_action_signals; // @[programmableCache.scala 434:41]
  assign compUnit_3_io_clear = _T_451 & actionReg_3_io_deq_valid; // @[programmableCache.scala 381:30]
  assign compUnit_3_io_op1_valid = compUnitInput1_3_io_out_valid; // @[programmableCache.scala 425:28]
  assign compUnit_3_io_op1_bits = compUnitInput1_3_io_out_bits; // @[programmableCache.scala 425:28]
  assign compUnit_3_io_op2_valid = compUnitInput2_3_io_out_valid; // @[programmableCache.scala 432:28]
  assign compUnit_3_io_op2_bits = compUnitInput2_3_io_out_bits; // @[programmableCache.scala 432:28]
  assign compUnit_4_clock = clock;
  assign compUnit_4_reset = reset;
  assign compUnit_4_io_instruction_valid = _T_512 & actionReg_4_io_deq_valid; // @[programmableCache.scala 435:42]
  assign compUnit_4_io_instruction_bits = actionReg_4_io_deq_bits_action_signals; // @[programmableCache.scala 434:41]
  assign compUnit_4_io_clear = _T_508 & actionReg_4_io_deq_valid; // @[programmableCache.scala 381:30]
  assign compUnit_4_io_op1_valid = compUnitInput1_4_io_out_valid; // @[programmableCache.scala 425:28]
  assign compUnit_4_io_op1_bits = compUnitInput1_4_io_out_bits; // @[programmableCache.scala 425:28]
  assign compUnit_4_io_op2_valid = compUnitInput2_4_io_out_valid; // @[programmableCache.scala 432:28]
  assign compUnit_4_io_op2_bits = compUnitInput2_4_io_out_bits; // @[programmableCache.scala 432:28]
  assign compUnit_5_clock = clock;
  assign compUnit_5_reset = reset;
  assign compUnit_5_io_instruction_valid = _T_569 & actionReg_5_io_deq_valid; // @[programmableCache.scala 435:42]
  assign compUnit_5_io_instruction_bits = actionReg_5_io_deq_bits_action_signals; // @[programmableCache.scala 434:41]
  assign compUnit_5_io_clear = _T_565 & actionReg_5_io_deq_valid; // @[programmableCache.scala 381:30]
  assign compUnit_5_io_op1_valid = compUnitInput1_5_io_out_valid; // @[programmableCache.scala 425:28]
  assign compUnit_5_io_op1_bits = compUnitInput1_5_io_out_bits; // @[programmableCache.scala 425:28]
  assign compUnit_5_io_op2_valid = compUnitInput2_5_io_out_valid; // @[programmableCache.scala 432:28]
  assign compUnit_5_io_op2_bits = compUnitInput2_5_io_out_bits; // @[programmableCache.scala 432:28]
  assign compUnit_6_clock = clock;
  assign compUnit_6_reset = reset;
  assign compUnit_6_io_instruction_valid = _T_626 & actionReg_6_io_deq_valid; // @[programmableCache.scala 435:42]
  assign compUnit_6_io_instruction_bits = actionReg_6_io_deq_bits_action_signals; // @[programmableCache.scala 434:41]
  assign compUnit_6_io_clear = _T_622 & actionReg_6_io_deq_valid; // @[programmableCache.scala 381:30]
  assign compUnit_6_io_op1_valid = compUnitInput1_6_io_out_valid; // @[programmableCache.scala 425:28]
  assign compUnit_6_io_op1_bits = compUnitInput1_6_io_out_bits; // @[programmableCache.scala 425:28]
  assign compUnit_6_io_op2_valid = compUnitInput2_6_io_out_valid; // @[programmableCache.scala 432:28]
  assign compUnit_6_io_op2_bits = compUnitInput2_6_io_out_bits; // @[programmableCache.scala 432:28]
  assign compUnit_7_clock = clock;
  assign compUnit_7_reset = reset;
  assign compUnit_7_io_instruction_valid = _T_683 & actionReg_7_io_deq_valid; // @[programmableCache.scala 435:42]
  assign compUnit_7_io_instruction_bits = actionReg_7_io_deq_bits_action_signals; // @[programmableCache.scala 434:41]
  assign compUnit_7_io_clear = _T_679 & actionReg_7_io_deq_valid; // @[programmableCache.scala 381:30]
  assign compUnit_7_io_op1_valid = compUnitInput1_7_io_out_valid; // @[programmableCache.scala 425:28]
  assign compUnit_7_io_op1_bits = compUnitInput1_7_io_out_bits; // @[programmableCache.scala 425:28]
  assign compUnit_7_io_op2_valid = compUnitInput2_7_io_out_valid; // @[programmableCache.scala 432:28]
  assign compUnit_7_io_op2_bits = compUnitInput2_7_io_out_bits; // @[programmableCache.scala 432:28]
  assign compUnitInput1_0_io_in_hardCoded = 64'h0;
  assign compUnitInput1_0_io_in_data = 64'h0;
  assign compUnitInput1_0_io_in_tbe = {{32'd0}, actionReg_0_io_deq_bits_addr}; // @[programmableCache.scala 422:38]
  assign compUnitInput1_0_io_in_select = {{1'd0}, actionReg_0_io_deq_bits_action_actionType[0]}; // @[programmableCache.scala 424:40]
  assign compUnitInput1_1_io_in_hardCoded = 64'h0;
  assign compUnitInput1_1_io_in_data = 64'h0;
  assign compUnitInput1_1_io_in_tbe = {{32'd0}, actionReg_1_io_deq_bits_addr}; // @[programmableCache.scala 422:38]
  assign compUnitInput1_1_io_in_select = {{1'd0}, actionReg_1_io_deq_bits_action_actionType[0]}; // @[programmableCache.scala 424:40]
  assign compUnitInput1_2_io_in_hardCoded = 64'h0;
  assign compUnitInput1_2_io_in_data = 64'h0;
  assign compUnitInput1_2_io_in_tbe = {{32'd0}, actionReg_2_io_deq_bits_addr}; // @[programmableCache.scala 422:38]
  assign compUnitInput1_2_io_in_select = {{1'd0}, actionReg_2_io_deq_bits_action_actionType[0]}; // @[programmableCache.scala 424:40]
  assign compUnitInput1_3_io_in_hardCoded = 64'h0;
  assign compUnitInput1_3_io_in_data = 64'h0;
  assign compUnitInput1_3_io_in_tbe = {{32'd0}, actionReg_3_io_deq_bits_addr}; // @[programmableCache.scala 422:38]
  assign compUnitInput1_3_io_in_select = {{1'd0}, actionReg_3_io_deq_bits_action_actionType[0]}; // @[programmableCache.scala 424:40]
  assign compUnitInput1_4_io_in_hardCoded = 64'h0;
  assign compUnitInput1_4_io_in_data = 64'h0;
  assign compUnitInput1_4_io_in_tbe = {{32'd0}, actionReg_4_io_deq_bits_addr}; // @[programmableCache.scala 422:38]
  assign compUnitInput1_4_io_in_select = {{1'd0}, actionReg_4_io_deq_bits_action_actionType[0]}; // @[programmableCache.scala 424:40]
  assign compUnitInput1_5_io_in_hardCoded = 64'h0;
  assign compUnitInput1_5_io_in_data = 64'h0;
  assign compUnitInput1_5_io_in_tbe = {{32'd0}, actionReg_5_io_deq_bits_addr}; // @[programmableCache.scala 422:38]
  assign compUnitInput1_5_io_in_select = {{1'd0}, actionReg_5_io_deq_bits_action_actionType[0]}; // @[programmableCache.scala 424:40]
  assign compUnitInput1_6_io_in_hardCoded = 64'h0;
  assign compUnitInput1_6_io_in_data = 64'h0;
  assign compUnitInput1_6_io_in_tbe = {{32'd0}, actionReg_6_io_deq_bits_addr}; // @[programmableCache.scala 422:38]
  assign compUnitInput1_6_io_in_select = {{1'd0}, actionReg_6_io_deq_bits_action_actionType[0]}; // @[programmableCache.scala 424:40]
  assign compUnitInput1_7_io_in_hardCoded = 64'h0;
  assign compUnitInput1_7_io_in_data = 64'h0;
  assign compUnitInput1_7_io_in_tbe = {{32'd0}, actionReg_7_io_deq_bits_addr}; // @[programmableCache.scala 422:38]
  assign compUnitInput1_7_io_in_select = {{1'd0}, actionReg_7_io_deq_bits_action_actionType[0]}; // @[programmableCache.scala 424:40]
  assign compUnitInput2_0_io_in_hardCoded = {{48'd0}, actionReg_0_io_deq_bits_action_signals[27:12]}; // @[programmableCache.scala 430:43]
  assign compUnitInput2_0_io_in_data = actionReg_0_io_deq_bits_data; // @[programmableCache.scala 428:38]
  assign compUnitInput2_0_io_in_tbe = {{32'd0}, actionReg_0_io_deq_bits_tbeFields_0}; // @[programmableCache.scala 429:38]
  assign compUnitInput2_0_io_in_select = actionReg_0_io_deq_bits_action_actionType[2:1]; // @[programmableCache.scala 431:40]
  assign compUnitInput2_1_io_in_hardCoded = {{48'd0}, actionReg_1_io_deq_bits_action_signals[27:12]}; // @[programmableCache.scala 430:43]
  assign compUnitInput2_1_io_in_data = actionReg_1_io_deq_bits_data; // @[programmableCache.scala 428:38]
  assign compUnitInput2_1_io_in_tbe = {{32'd0}, actionReg_1_io_deq_bits_tbeFields_0}; // @[programmableCache.scala 429:38]
  assign compUnitInput2_1_io_in_select = actionReg_1_io_deq_bits_action_actionType[2:1]; // @[programmableCache.scala 431:40]
  assign compUnitInput2_2_io_in_hardCoded = {{48'd0}, actionReg_2_io_deq_bits_action_signals[27:12]}; // @[programmableCache.scala 430:43]
  assign compUnitInput2_2_io_in_data = actionReg_2_io_deq_bits_data; // @[programmableCache.scala 428:38]
  assign compUnitInput2_2_io_in_tbe = {{32'd0}, actionReg_2_io_deq_bits_tbeFields_0}; // @[programmableCache.scala 429:38]
  assign compUnitInput2_2_io_in_select = actionReg_2_io_deq_bits_action_actionType[2:1]; // @[programmableCache.scala 431:40]
  assign compUnitInput2_3_io_in_hardCoded = {{48'd0}, actionReg_3_io_deq_bits_action_signals[27:12]}; // @[programmableCache.scala 430:43]
  assign compUnitInput2_3_io_in_data = actionReg_3_io_deq_bits_data; // @[programmableCache.scala 428:38]
  assign compUnitInput2_3_io_in_tbe = {{32'd0}, actionReg_3_io_deq_bits_tbeFields_0}; // @[programmableCache.scala 429:38]
  assign compUnitInput2_3_io_in_select = actionReg_3_io_deq_bits_action_actionType[2:1]; // @[programmableCache.scala 431:40]
  assign compUnitInput2_4_io_in_hardCoded = {{48'd0}, actionReg_4_io_deq_bits_action_signals[27:12]}; // @[programmableCache.scala 430:43]
  assign compUnitInput2_4_io_in_data = actionReg_4_io_deq_bits_data; // @[programmableCache.scala 428:38]
  assign compUnitInput2_4_io_in_tbe = {{32'd0}, actionReg_4_io_deq_bits_tbeFields_0}; // @[programmableCache.scala 429:38]
  assign compUnitInput2_4_io_in_select = actionReg_4_io_deq_bits_action_actionType[2:1]; // @[programmableCache.scala 431:40]
  assign compUnitInput2_5_io_in_hardCoded = {{48'd0}, actionReg_5_io_deq_bits_action_signals[27:12]}; // @[programmableCache.scala 430:43]
  assign compUnitInput2_5_io_in_data = actionReg_5_io_deq_bits_data; // @[programmableCache.scala 428:38]
  assign compUnitInput2_5_io_in_tbe = {{32'd0}, actionReg_5_io_deq_bits_tbeFields_0}; // @[programmableCache.scala 429:38]
  assign compUnitInput2_5_io_in_select = actionReg_5_io_deq_bits_action_actionType[2:1]; // @[programmableCache.scala 431:40]
  assign compUnitInput2_6_io_in_hardCoded = {{48'd0}, actionReg_6_io_deq_bits_action_signals[27:12]}; // @[programmableCache.scala 430:43]
  assign compUnitInput2_6_io_in_data = actionReg_6_io_deq_bits_data; // @[programmableCache.scala 428:38]
  assign compUnitInput2_6_io_in_tbe = {{32'd0}, actionReg_6_io_deq_bits_tbeFields_0}; // @[programmableCache.scala 429:38]
  assign compUnitInput2_6_io_in_select = actionReg_6_io_deq_bits_action_actionType[2:1]; // @[programmableCache.scala 431:40]
  assign compUnitInput2_7_io_in_hardCoded = {{48'd0}, actionReg_7_io_deq_bits_action_signals[27:12]}; // @[programmableCache.scala 430:43]
  assign compUnitInput2_7_io_in_data = actionReg_7_io_deq_bits_data; // @[programmableCache.scala 428:38]
  assign compUnitInput2_7_io_in_tbe = {{32'd0}, actionReg_7_io_deq_bits_tbeFields_0}; // @[programmableCache.scala 429:38]
  assign compUnitInput2_7_io_in_select = actionReg_7_io_deq_bits_action_actionType[2:1]; // @[programmableCache.scala 431:40]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  instUsed = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  replStateReg_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  replStateReg_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  wayInputCache = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  tbeFields_0 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  _T_270 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  inputToPC_addr = _RAND_6[31:0];
  _RAND_7 = {2{`RANDOM}};
  inputToPC_data = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  _T_783 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  _T_785 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  _T_786 = _RAND_10[31:0];
  _RAND_11 = {2{`RANDOM}};
  _T_787 = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  _T_790 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  _T_798 = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      instUsed <= 1'h0;
    end else begin
      instUsed <= _T_170;
    end
    if (reset) begin
      replStateReg_0 <= 1'h0;
    end else if (missLD) begin
      if (~addrReplacer[0]) begin
        replStateReg_0 <= _T_261[1];
      end
    end
    if (reset) begin
      replStateReg_1 <= 1'h0;
    end else if (missLD) begin
      if (addrReplacer[0]) begin
        replStateReg_1 <= _T_261[1];
      end
    end
    if (reset) begin
      wayInputCache <= 3'h2;
    end else if (getState) begin
      if (_T_263) begin
        wayInputCache <= {{1'd0}, probeWay_io_deq_bits};
      end else begin
        wayInputCache <= tbeWay;
      end
    end
    if (reset) begin
      tbeFields_0 <= 32'h0;
    end else if (getState) begin
      tbeFields_0 <= input__io_deq_bits_tbeOut_fields_0;
    end
    if (reset) begin
      _T_270 <= 2'h2;
    end else if (getState) begin
      _T_270 <= {{1'd0}, replacerWayWire};
    end
    if (reset) begin
      inputToPC_addr <= 32'h0;
    end else if (getState) begin
      inputToPC_addr <= input__io_deq_bits_inst_addr;
    end
    if (reset) begin
      inputToPC_data <= 64'h0;
    end else if (getState) begin
      inputToPC_data <= input__io_deq_bits_inst_data;
    end
    _T_783 <= cache_io_bipassLD_in_bits_addr;
    _T_785 <= inputArbiter_io_chosen;
    _T_786 <= inputArbiter_io_out_bits_addr;
    _T_787 <= inputArbiter_io_out_bits_data;
    _T_790 <= inputArbiter_io_chosen;
    _T_798 <= tbe_io_isFull;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_784 & _T_789) begin
          $fwrite(32'h80000002,"Cache: %d req from %d Addr: %d Data: %d\n",1'h0,_T_785,_T_786,_T_787); // @[programmableCache.scala 531:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1543 & _T_789) begin
          $fwrite(32'h80000002,"Cache: %d ",1'h0); // @[programmableCache.scala 533:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1545 & _T_789) begin
          $fwrite(32'h80000002," Load hit for addr %d\n",input__io_deq_bits_inst_addr); // @[programmableCache.scala 535:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1549 & _T_789) begin
          $fwrite(32'h80000002,"addr %d is locked\n",input__io_deq_bits_inst_addr); // @[programmableCache.scala 537:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1555 & _T_789) begin
          $fwrite(32'h80000002,"TBE is full addr %d\n",input__io_deq_bits_inst_addr); // @[programmableCache.scala 539:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1563 & _T_789) begin
          $fwrite(32'h80000002,"Hit (store probably) for addr %d\n",input__io_deq_bits_inst_addr); // @[programmableCache.scala 541:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1572 & _T_789) begin
          $fwrite(32'h80000002,"miss for addr %d\n",input__io_deq_bits_inst_addr); // @[programmableCache.scala 543:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (getState & _T_789) begin
          $fwrite(32'h80000002,"Event %d Addr: %d Data: %d\n",input__io_deq_bits_inst_event,input__io_deq_bits_inst_addr,input__io_deq_bits_inst_data); // @[programmableCache.scala 549:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CacheNode(
  input         clock,
  input         reset,
  output        io_in_cpu_ready,
  input         io_in_cpu_valid,
  input  [31:0] io_in_cpu_bits_addr,
  input  [7:0]  io_in_cpu_bits_inst,
  input  [63:0] io_in_cpu_bits_data,
  output        io_in_network_ready,
  input         io_in_network_valid,
  input  [31:0] io_in_network_bits_addr,
  input  [7:0]  io_in_network_bits_inst,
  input  [63:0] io_in_network_bits_data,
  input  [1:0]  io_in_network_bits_msgType,
  output        io_out_network_valid,
  output [31:0] io_out_network_bits_addr,
  output [7:0]  io_out_network_bits_inst,
  output [63:0] io_out_network_bits_data,
  output        io_out_cpu_valid,
  output [31:0] io_out_cpu_bits_addr,
  output        _T_814,
  output        _T_808,
  output        _T_819,
  output        hitLD,
  output        missLD,
  output        _T_811
);
  wire  cache_clock; // @[cacheNode.scala 33:21]
  wire  cache_reset; // @[cacheNode.scala 33:21]
  wire  cache_io_in_cpu_ready; // @[cacheNode.scala 33:21]
  wire  cache_io_in_cpu_valid; // @[cacheNode.scala 33:21]
  wire [1:0] cache_io_in_cpu_bits_event; // @[cacheNode.scala 33:21]
  wire [31:0] cache_io_in_cpu_bits_addr; // @[cacheNode.scala 33:21]
  wire [63:0] cache_io_in_cpu_bits_data; // @[cacheNode.scala 33:21]
  wire  cache_io_in_memCtrl_ready; // @[cacheNode.scala 33:21]
  wire  cache_io_in_memCtrl_valid; // @[cacheNode.scala 33:21]
  wire [1:0] cache_io_in_memCtrl_bits_event; // @[cacheNode.scala 33:21]
  wire [31:0] cache_io_in_memCtrl_bits_addr; // @[cacheNode.scala 33:21]
  wire [63:0] cache_io_in_memCtrl_bits_data; // @[cacheNode.scala 33:21]
  wire  cache_io_in_otherNodes_ready; // @[cacheNode.scala 33:21]
  wire  cache_io_in_otherNodes_valid; // @[cacheNode.scala 33:21]
  wire [1:0] cache_io_in_otherNodes_bits_event; // @[cacheNode.scala 33:21]
  wire [31:0] cache_io_in_otherNodes_bits_addr; // @[cacheNode.scala 33:21]
  wire [63:0] cache_io_in_otherNodes_bits_data; // @[cacheNode.scala 33:21]
  wire  cache_io_out_req_valid; // @[cacheNode.scala 33:21]
  wire [31:0] cache_io_out_req_bits_req_addr; // @[cacheNode.scala 33:21]
  wire [7:0] cache_io_out_req_bits_req_inst; // @[cacheNode.scala 33:21]
  wire [63:0] cache_io_out_req_bits_req_data; // @[cacheNode.scala 33:21]
  wire  cache_io_out_resp_valid; // @[cacheNode.scala 33:21]
  wire [31:0] cache_io_out_resp_bits_addr; // @[cacheNode.scala 33:21]
  wire  cache__T_814_0; // @[cacheNode.scala 33:21]
  wire  cache__T_808_0; // @[cacheNode.scala 33:21]
  wire  cache__T_819_0; // @[cacheNode.scala 33:21]
  wire  cache_hitLD_0; // @[cacheNode.scala 33:21]
  wire  cache_missLD_0; // @[cacheNode.scala 33:21]
  wire  cache__T_811_0; // @[cacheNode.scala 33:21]
  wire  cpuQueue_clock; // @[cacheNode.scala 34:24]
  wire  cpuQueue_reset; // @[cacheNode.scala 34:24]
  wire  cpuQueue_io_enq_ready; // @[cacheNode.scala 34:24]
  wire  cpuQueue_io_enq_valid; // @[cacheNode.scala 34:24]
  wire [31:0] cpuQueue_io_enq_bits_addr; // @[cacheNode.scala 34:24]
  wire [7:0] cpuQueue_io_enq_bits_inst; // @[cacheNode.scala 34:24]
  wire [63:0] cpuQueue_io_enq_bits_data; // @[cacheNode.scala 34:24]
  wire  cpuQueue_io_deq_ready; // @[cacheNode.scala 34:24]
  wire  cpuQueue_io_deq_valid; // @[cacheNode.scala 34:24]
  wire [31:0] cpuQueue_io_deq_bits_addr; // @[cacheNode.scala 34:24]
  wire [7:0] cpuQueue_io_deq_bits_inst; // @[cacheNode.scala 34:24]
  wire [63:0] cpuQueue_io_deq_bits_data; // @[cacheNode.scala 34:24]
  wire  memCtrlQueue_clock; // @[cacheNode.scala 35:28]
  wire  memCtrlQueue_reset; // @[cacheNode.scala 35:28]
  wire  memCtrlQueue_io_enq_ready; // @[cacheNode.scala 35:28]
  wire  memCtrlQueue_io_enq_valid; // @[cacheNode.scala 35:28]
  wire [31:0] memCtrlQueue_io_enq_bits_addr; // @[cacheNode.scala 35:28]
  wire [7:0] memCtrlQueue_io_enq_bits_inst; // @[cacheNode.scala 35:28]
  wire [63:0] memCtrlQueue_io_enq_bits_data; // @[cacheNode.scala 35:28]
  wire  memCtrlQueue_io_deq_ready; // @[cacheNode.scala 35:28]
  wire  memCtrlQueue_io_deq_valid; // @[cacheNode.scala 35:28]
  wire [31:0] memCtrlQueue_io_deq_bits_addr; // @[cacheNode.scala 35:28]
  wire [7:0] memCtrlQueue_io_deq_bits_inst; // @[cacheNode.scala 35:28]
  wire [63:0] memCtrlQueue_io_deq_bits_data; // @[cacheNode.scala 35:28]
  wire  otherNodesQueue_clock; // @[cacheNode.scala 36:31]
  wire  otherNodesQueue_reset; // @[cacheNode.scala 36:31]
  wire  otherNodesQueue_io_enq_ready; // @[cacheNode.scala 36:31]
  wire  otherNodesQueue_io_enq_valid; // @[cacheNode.scala 36:31]
  wire [31:0] otherNodesQueue_io_enq_bits_addr; // @[cacheNode.scala 36:31]
  wire [7:0] otherNodesQueue_io_enq_bits_inst; // @[cacheNode.scala 36:31]
  wire [63:0] otherNodesQueue_io_enq_bits_data; // @[cacheNode.scala 36:31]
  wire  otherNodesQueue_io_deq_ready; // @[cacheNode.scala 36:31]
  wire  otherNodesQueue_io_deq_valid; // @[cacheNode.scala 36:31]
  wire [31:0] otherNodesQueue_io_deq_bits_addr; // @[cacheNode.scala 36:31]
  wire [7:0] otherNodesQueue_io_deq_bits_inst; // @[cacheNode.scala 36:31]
  wire [63:0] otherNodesQueue_io_deq_bits_data; // @[cacheNode.scala 36:31]
  wire  _T_1 = io_in_network_ready & io_in_network_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_in_network_bits_msgType == 2'h0; // @[cacheNode.scala 54:37]
  wire  _T_3 = io_in_network_bits_msgType == 2'h1; // @[cacheNode.scala 56:43]
  wire  _GEN_2 = _T_2 ? 1'h0 : _T_3; // @[cacheNode.scala 54:45]
  programmableCache cache ( // @[cacheNode.scala 33:21]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_in_cpu_ready(cache_io_in_cpu_ready),
    .io_in_cpu_valid(cache_io_in_cpu_valid),
    .io_in_cpu_bits_event(cache_io_in_cpu_bits_event),
    .io_in_cpu_bits_addr(cache_io_in_cpu_bits_addr),
    .io_in_cpu_bits_data(cache_io_in_cpu_bits_data),
    .io_in_memCtrl_ready(cache_io_in_memCtrl_ready),
    .io_in_memCtrl_valid(cache_io_in_memCtrl_valid),
    .io_in_memCtrl_bits_event(cache_io_in_memCtrl_bits_event),
    .io_in_memCtrl_bits_addr(cache_io_in_memCtrl_bits_addr),
    .io_in_memCtrl_bits_data(cache_io_in_memCtrl_bits_data),
    .io_in_otherNodes_ready(cache_io_in_otherNodes_ready),
    .io_in_otherNodes_valid(cache_io_in_otherNodes_valid),
    .io_in_otherNodes_bits_event(cache_io_in_otherNodes_bits_event),
    .io_in_otherNodes_bits_addr(cache_io_in_otherNodes_bits_addr),
    .io_in_otherNodes_bits_data(cache_io_in_otherNodes_bits_data),
    .io_out_req_valid(cache_io_out_req_valid),
    .io_out_req_bits_req_addr(cache_io_out_req_bits_req_addr),
    .io_out_req_bits_req_inst(cache_io_out_req_bits_req_inst),
    .io_out_req_bits_req_data(cache_io_out_req_bits_req_data),
    .io_out_resp_valid(cache_io_out_resp_valid),
    .io_out_resp_bits_addr(cache_io_out_resp_bits_addr),
    ._T_814_0(cache__T_814_0),
    ._T_808_0(cache__T_808_0),
    ._T_819_0(cache__T_819_0),
    .hitLD_0(cache_hitLD_0),
    .missLD_0(cache_missLD_0),
    ._T_811_0(cache__T_811_0)
  );
  Queue_17 cpuQueue ( // @[cacheNode.scala 34:24]
    .clock(cpuQueue_clock),
    .reset(cpuQueue_reset),
    .io_enq_ready(cpuQueue_io_enq_ready),
    .io_enq_valid(cpuQueue_io_enq_valid),
    .io_enq_bits_addr(cpuQueue_io_enq_bits_addr),
    .io_enq_bits_inst(cpuQueue_io_enq_bits_inst),
    .io_enq_bits_data(cpuQueue_io_enq_bits_data),
    .io_deq_ready(cpuQueue_io_deq_ready),
    .io_deq_valid(cpuQueue_io_deq_valid),
    .io_deq_bits_addr(cpuQueue_io_deq_bits_addr),
    .io_deq_bits_inst(cpuQueue_io_deq_bits_inst),
    .io_deq_bits_data(cpuQueue_io_deq_bits_data)
  );
  Queue_17 memCtrlQueue ( // @[cacheNode.scala 35:28]
    .clock(memCtrlQueue_clock),
    .reset(memCtrlQueue_reset),
    .io_enq_ready(memCtrlQueue_io_enq_ready),
    .io_enq_valid(memCtrlQueue_io_enq_valid),
    .io_enq_bits_addr(memCtrlQueue_io_enq_bits_addr),
    .io_enq_bits_inst(memCtrlQueue_io_enq_bits_inst),
    .io_enq_bits_data(memCtrlQueue_io_enq_bits_data),
    .io_deq_ready(memCtrlQueue_io_deq_ready),
    .io_deq_valid(memCtrlQueue_io_deq_valid),
    .io_deq_bits_addr(memCtrlQueue_io_deq_bits_addr),
    .io_deq_bits_inst(memCtrlQueue_io_deq_bits_inst),
    .io_deq_bits_data(memCtrlQueue_io_deq_bits_data)
  );
  Queue_17 otherNodesQueue ( // @[cacheNode.scala 36:31]
    .clock(otherNodesQueue_clock),
    .reset(otherNodesQueue_reset),
    .io_enq_ready(otherNodesQueue_io_enq_ready),
    .io_enq_valid(otherNodesQueue_io_enq_valid),
    .io_enq_bits_addr(otherNodesQueue_io_enq_bits_addr),
    .io_enq_bits_inst(otherNodesQueue_io_enq_bits_inst),
    .io_enq_bits_data(otherNodesQueue_io_enq_bits_data),
    .io_deq_ready(otherNodesQueue_io_deq_ready),
    .io_deq_valid(otherNodesQueue_io_deq_valid),
    .io_deq_bits_addr(otherNodesQueue_io_deq_bits_addr),
    .io_deq_bits_inst(otherNodesQueue_io_deq_bits_inst),
    .io_deq_bits_data(otherNodesQueue_io_deq_bits_data)
  );
  assign io_in_cpu_ready = cpuQueue_io_enq_ready; // @[cacheNode.scala 38:19]
  assign io_in_network_ready = memCtrlQueue_io_enq_ready & otherNodesQueue_io_enq_ready; // @[cacheNode.scala 47:23]
  assign io_out_network_valid = cache_io_out_req_valid; // @[cacheNode.scala 81:24]
  assign io_out_network_bits_addr = cache_io_out_req_bits_req_addr; // @[cacheNode.scala 86:28]
  assign io_out_network_bits_inst = cache_io_out_req_bits_req_inst; // @[cacheNode.scala 84:27]
  assign io_out_network_bits_data = cache_io_out_req_bits_req_data; // @[cacheNode.scala 85:28]
  assign io_out_cpu_valid = cache_io_out_resp_valid; // @[cacheNode.scala 92:20]
  assign io_out_cpu_bits_addr = cache_io_out_resp_bits_addr; // @[cacheNode.scala 90:24]
  assign _T_814 = cache__T_814_0;
  assign _T_808 = cache__T_808_0;
  assign _T_819 = cache__T_819_0;
  assign hitLD = cache_hitLD_0;
  assign missLD = cache_missLD_0;
  assign _T_811 = cache__T_811_0;
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_in_cpu_valid = cpuQueue_io_deq_valid; // @[cacheNode.scala 64:30]
  assign cache_io_in_cpu_bits_event = cpuQueue_io_deq_bits_inst[1:0]; // @[cacheNode.scala 61:30]
  assign cache_io_in_cpu_bits_addr = cpuQueue_io_deq_bits_addr; // @[cacheNode.scala 62:30]
  assign cache_io_in_cpu_bits_data = cpuQueue_io_deq_bits_data; // @[cacheNode.scala 63:30]
  assign cache_io_in_memCtrl_valid = memCtrlQueue_io_deq_valid; // @[cacheNode.scala 70:34]
  assign cache_io_in_memCtrl_bits_event = memCtrlQueue_io_deq_bits_inst[1:0]; // @[cacheNode.scala 67:34]
  assign cache_io_in_memCtrl_bits_addr = memCtrlQueue_io_deq_bits_addr; // @[cacheNode.scala 68:34]
  assign cache_io_in_memCtrl_bits_data = memCtrlQueue_io_deq_bits_data; // @[cacheNode.scala 69:34]
  assign cache_io_in_otherNodes_valid = otherNodesQueue_io_deq_valid; // @[cacheNode.scala 76:37]
  assign cache_io_in_otherNodes_bits_event = otherNodesQueue_io_deq_bits_inst[1:0]; // @[cacheNode.scala 73:37]
  assign cache_io_in_otherNodes_bits_addr = otherNodesQueue_io_deq_bits_addr; // @[cacheNode.scala 74:37]
  assign cache_io_in_otherNodes_bits_data = otherNodesQueue_io_deq_bits_data; // @[cacheNode.scala 75:37]
  assign cpuQueue_clock = clock;
  assign cpuQueue_reset = reset;
  assign cpuQueue_io_enq_valid = io_in_cpu_valid; // @[cacheNode.scala 38:19]
  assign cpuQueue_io_enq_bits_addr = io_in_cpu_bits_addr; // @[cacheNode.scala 38:19]
  assign cpuQueue_io_enq_bits_inst = io_in_cpu_bits_inst; // @[cacheNode.scala 38:19]
  assign cpuQueue_io_enq_bits_data = io_in_cpu_bits_data; // @[cacheNode.scala 38:19]
  assign cpuQueue_io_deq_ready = cache_io_in_cpu_ready; // @[cacheNode.scala 65:25]
  assign memCtrlQueue_clock = clock;
  assign memCtrlQueue_reset = reset;
  assign memCtrlQueue_io_enq_valid = _T_1 & _T_2; // @[cacheNode.scala 49:29 cacheNode.scala 55:33]
  assign memCtrlQueue_io_enq_bits_addr = io_in_network_bits_addr; // @[cacheNode.scala 39:33]
  assign memCtrlQueue_io_enq_bits_inst = io_in_network_bits_inst; // @[cacheNode.scala 41:33]
  assign memCtrlQueue_io_enq_bits_data = io_in_network_bits_data; // @[cacheNode.scala 40:33]
  assign memCtrlQueue_io_deq_ready = cache_io_in_memCtrl_ready; // @[cacheNode.scala 71:29]
  assign otherNodesQueue_clock = clock;
  assign otherNodesQueue_reset = reset;
  assign otherNodesQueue_io_enq_valid = _T_1 & _GEN_2; // @[cacheNode.scala 50:32 cacheNode.scala 57:36]
  assign otherNodesQueue_io_enq_bits_addr = io_in_network_bits_addr; // @[cacheNode.scala 43:36]
  assign otherNodesQueue_io_enq_bits_inst = io_in_network_bits_inst; // @[cacheNode.scala 45:36]
  assign otherNodesQueue_io_enq_bits_data = io_in_network_bits_data; // @[cacheNode.scala 44:36]
  assign otherNodesQueue_io_deq_ready = cache_io_in_otherNodes_ready; // @[cacheNode.scala 77:32]
endmodule
module Bore(
  input         clock,
  input         reset,
  output [31:0] io_events_0,
  output [31:0] io_events_1,
  output [31:0] io_events_2,
  output [31:0] io_events_3,
  output [31:0] io_events_4,
  output [31:0] io_events_5,
  input         memCtrlReq_0,
  input         instCount_0,
  input         ldReq_0,
  input         hitLD_0,
  input         missLD_0,
  input         cpuReq_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [23:0] _T_1; // @[Counter.scala 29:33]
  wire  _T_3 = _T_1 == 24'h98967f; // @[Counter.scala 38:24]
  wire [23:0] _T_5 = _T_1 + 24'h1; // @[Counter.scala 39:22]
  reg [23:0] _T_6; // @[Counter.scala 29:33]
  wire  _T_8 = _T_6 == 24'h98967f; // @[Counter.scala 38:24]
  wire [23:0] _T_10 = _T_6 + 24'h1; // @[Counter.scala 39:22]
  reg [23:0] _T_11; // @[Counter.scala 29:33]
  wire  _T_13 = _T_11 == 24'h98967f; // @[Counter.scala 38:24]
  wire [23:0] _T_15 = _T_11 + 24'h1; // @[Counter.scala 39:22]
  reg [23:0] _T_16; // @[Counter.scala 29:33]
  wire  _T_18 = _T_16 == 24'h98967f; // @[Counter.scala 38:24]
  wire [23:0] _T_20 = _T_16 + 24'h1; // @[Counter.scala 39:22]
  reg [23:0] _T_21; // @[Counter.scala 29:33]
  wire  _T_23 = _T_21 == 24'h98967f; // @[Counter.scala 38:24]
  wire [23:0] _T_25 = _T_21 + 24'h1; // @[Counter.scala 39:22]
  reg [23:0] _T_26; // @[Counter.scala 29:33]
  wire  _T_28 = _T_26 == 24'h98967f; // @[Counter.scala 38:24]
  wire [23:0] _T_30 = _T_26 + 24'h1; // @[Counter.scala 39:22]
  assign io_events_0 = {{8'd0}, _T_1}; // @[memGenTopLevel.scala 40:15]
  assign io_events_1 = {{8'd0}, _T_6}; // @[memGenTopLevel.scala 40:15]
  assign io_events_2 = {{8'd0}, _T_11}; // @[memGenTopLevel.scala 40:15]
  assign io_events_3 = {{8'd0}, _T_16}; // @[memGenTopLevel.scala 40:15]
  assign io_events_4 = {{8'd0}, _T_21}; // @[memGenTopLevel.scala 40:15]
  assign io_events_5 = {{8'd0}, _T_26}; // @[memGenTopLevel.scala 40:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[23:0];
  _RAND_1 = {1{`RANDOM}};
  _T_6 = _RAND_1[23:0];
  _RAND_2 = {1{`RANDOM}};
  _T_11 = _RAND_2[23:0];
  _RAND_3 = {1{`RANDOM}};
  _T_16 = _RAND_3[23:0];
  _RAND_4 = {1{`RANDOM}};
  _T_21 = _RAND_4[23:0];
  _RAND_5 = {1{`RANDOM}};
  _T_26 = _RAND_5[23:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1 <= 24'h0;
    end else if (missLD_0) begin
      if (_T_3) begin
        _T_1 <= 24'h0;
      end else begin
        _T_1 <= _T_5;
      end
    end
    if (reset) begin
      _T_6 <= 24'h0;
    end else if (hitLD_0) begin
      if (_T_8) begin
        _T_6 <= 24'h0;
      end else begin
        _T_6 <= _T_10;
      end
    end
    if (reset) begin
      _T_11 <= 24'h0;
    end else if (instCount_0) begin
      if (_T_13) begin
        _T_11 <= 24'h0;
      end else begin
        _T_11 <= _T_15;
      end
    end
    if (reset) begin
      _T_16 <= 24'h0;
    end else if (cpuReq_0) begin
      if (_T_18) begin
        _T_16 <= 24'h0;
      end else begin
        _T_16 <= _T_20;
      end
    end
    if (reset) begin
      _T_21 <= 24'h0;
    end else if (memCtrlReq_0) begin
      if (_T_23) begin
        _T_21 <= 24'h0;
      end else begin
        _T_21 <= _T_25;
      end
    end
    if (reset) begin
      _T_26 <= 24'h0;
    end else if (ldReq_0) begin
      if (_T_28) begin
        _T_26 <= 24'h0;
      end else begin
        _T_26 <= _T_30;
      end
    end
  end
endmodule
module memGenTopLevel(
  input         clock,
  input         reset,
  output        io_instruction_0_ready,
  input         io_instruction_0_valid,
  input  [31:0] io_instruction_0_bits_addr,
  input  [7:0]  io_instruction_0_bits_inst,
  input  [63:0] io_instruction_0_bits_data,
  output        io_resp_0_valid,
  output [31:0] io_resp_0_bits_addr,
  output [31:0] io_events_bits_0,
  output [31:0] io_events_bits_1,
  output [31:0] io_events_bits_2,
  output [31:0] io_events_bits_3,
  output [31:0] io_events_bits_4,
  output [31:0] io_events_bits_5,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output        io_mem_b_ready,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [15:0] io_mem_ar_bits_len,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last
);
  wire  memCtrl_clock; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_reset; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_in_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_in_valid; // @[memGenTopLevel.scala 67:25]
  wire [31:0] memCtrl_io_in_bits_addr; // @[memGenTopLevel.scala 67:25]
  wire [7:0] memCtrl_io_in_bits_inst; // @[memGenTopLevel.scala 67:25]
  wire [63:0] memCtrl_io_in_bits_data; // @[memGenTopLevel.scala 67:25]
  wire [2:0] memCtrl_io_in_bits_src; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_aw_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_aw_valid; // @[memGenTopLevel.scala 67:25]
  wire [31:0] memCtrl_io_mem_aw_bits_addr; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_w_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_w_valid; // @[memGenTopLevel.scala 67:25]
  wire [63:0] memCtrl_io_mem_w_bits_data; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_b_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_ar_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_ar_valid; // @[memGenTopLevel.scala 67:25]
  wire [31:0] memCtrl_io_mem_ar_bits_addr; // @[memGenTopLevel.scala 67:25]
  wire [15:0] memCtrl_io_mem_ar_bits_len; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_r_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_r_valid; // @[memGenTopLevel.scala 67:25]
  wire [63:0] memCtrl_io_mem_r_bits_data; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_r_bits_last; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_out_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_out_valid; // @[memGenTopLevel.scala 67:25]
  wire [31:0] memCtrl_io_out_bits_addr; // @[memGenTopLevel.scala 67:25]
  wire [63:0] memCtrl_io_out_bits_data; // @[memGenTopLevel.scala 67:25]
  wire [2:0] memCtrl_io_out_bits_dst; // @[memGenTopLevel.scala 67:25]
  wire  memCtrlInputQueue_clock; // @[memGenTopLevel.scala 68:35]
  wire  memCtrlInputQueue_reset; // @[memGenTopLevel.scala 68:35]
  wire  memCtrlInputQueue_io_enq_ready; // @[memGenTopLevel.scala 68:35]
  wire  memCtrlInputQueue_io_enq_valid; // @[memGenTopLevel.scala 68:35]
  wire [31:0] memCtrlInputQueue_io_enq_bits_addr; // @[memGenTopLevel.scala 68:35]
  wire [7:0] memCtrlInputQueue_io_enq_bits_inst; // @[memGenTopLevel.scala 68:35]
  wire [63:0] memCtrlInputQueue_io_enq_bits_data; // @[memGenTopLevel.scala 68:35]
  wire [2:0] memCtrlInputQueue_io_enq_bits_src; // @[memGenTopLevel.scala 68:35]
  wire  memCtrlInputQueue_io_deq_ready; // @[memGenTopLevel.scala 68:35]
  wire  memCtrlInputQueue_io_deq_valid; // @[memGenTopLevel.scala 68:35]
  wire [31:0] memCtrlInputQueue_io_deq_bits_addr; // @[memGenTopLevel.scala 68:35]
  wire [7:0] memCtrlInputQueue_io_deq_bits_inst; // @[memGenTopLevel.scala 68:35]
  wire [63:0] memCtrlInputQueue_io_deq_bits_data; // @[memGenTopLevel.scala 68:35]
  wire [2:0] memCtrlInputQueue_io_deq_bits_src; // @[memGenTopLevel.scala 68:35]
  wire  routerNode_0_clock; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_reset; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_cacheIn_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_0_io_cacheIn_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_0_io_cacheIn_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_0_io_cacheIn_bits_data; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_cacheOut_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_cacheOut_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_0_io_cacheOut_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_0_io_cacheOut_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_0_io_cacheOut_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [1:0] routerNode_0_io_cacheOut_bits_msgType; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_in_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_in_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_0_io_in_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_0_io_in_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_0_io_in_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_0_io_in_bits_src; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_0_io_in_bits_dst; // @[memGenTopLevel.scala 70:28]
  wire [1:0] routerNode_0_io_in_bits_msgType; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_out_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_out_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_0_io_out_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_0_io_out_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_0_io_out_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_0_io_out_bits_src; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_0_io_out_bits_dst; // @[memGenTopLevel.scala 70:28]
  wire [1:0] routerNode_0_io_out_bits_msgType; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_clock; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_reset; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_cacheIn_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_cacheIn_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_1_io_cacheIn_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_1_io_cacheIn_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_1_io_cacheIn_bits_dst; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_cacheOut_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_cacheOut_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_1_io_cacheOut_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_1_io_cacheOut_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_1_io_cacheOut_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_1_io_cacheOut_bits_src; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_in_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_in_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_1_io_in_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_1_io_in_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_1_io_in_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_1_io_in_bits_src; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_1_io_in_bits_dst; // @[memGenTopLevel.scala 70:28]
  wire [1:0] routerNode_1_io_in_bits_msgType; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_out_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_out_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_1_io_out_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_1_io_out_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_1_io_out_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_1_io_out_bits_src; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_1_io_out_bits_dst; // @[memGenTopLevel.scala 70:28]
  wire [1:0] routerNode_1_io_out_bits_msgType; // @[memGenTopLevel.scala 70:28]
  wire  cacheNode_0_clock; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_reset; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_io_in_cpu_ready; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_io_in_cpu_valid; // @[memGenTopLevel.scala 74:28]
  wire [31:0] cacheNode_0_io_in_cpu_bits_addr; // @[memGenTopLevel.scala 74:28]
  wire [7:0] cacheNode_0_io_in_cpu_bits_inst; // @[memGenTopLevel.scala 74:28]
  wire [63:0] cacheNode_0_io_in_cpu_bits_data; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_io_in_network_ready; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_io_in_network_valid; // @[memGenTopLevel.scala 74:28]
  wire [31:0] cacheNode_0_io_in_network_bits_addr; // @[memGenTopLevel.scala 74:28]
  wire [7:0] cacheNode_0_io_in_network_bits_inst; // @[memGenTopLevel.scala 74:28]
  wire [63:0] cacheNode_0_io_in_network_bits_data; // @[memGenTopLevel.scala 74:28]
  wire [1:0] cacheNode_0_io_in_network_bits_msgType; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_io_out_network_valid; // @[memGenTopLevel.scala 74:28]
  wire [31:0] cacheNode_0_io_out_network_bits_addr; // @[memGenTopLevel.scala 74:28]
  wire [7:0] cacheNode_0_io_out_network_bits_inst; // @[memGenTopLevel.scala 74:28]
  wire [63:0] cacheNode_0_io_out_network_bits_data; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_io_out_cpu_valid; // @[memGenTopLevel.scala 74:28]
  wire [31:0] cacheNode_0_io_out_cpu_bits_addr; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0__T_814; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0__T_808; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0__T_819; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_hitLD; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_missLD; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0__T_811; // @[memGenTopLevel.scala 74:28]
  wire  bore_clock; // @[memGenTopLevel.scala 78:22]
  wire  bore_reset; // @[memGenTopLevel.scala 78:22]
  wire [31:0] bore_io_events_0; // @[memGenTopLevel.scala 78:22]
  wire [31:0] bore_io_events_1; // @[memGenTopLevel.scala 78:22]
  wire [31:0] bore_io_events_2; // @[memGenTopLevel.scala 78:22]
  wire [31:0] bore_io_events_3; // @[memGenTopLevel.scala 78:22]
  wire [31:0] bore_io_events_4; // @[memGenTopLevel.scala 78:22]
  wire [31:0] bore_io_events_5; // @[memGenTopLevel.scala 78:22]
  wire  bore_memCtrlReq_0; // @[memGenTopLevel.scala 78:22]
  wire  bore_instCount_0; // @[memGenTopLevel.scala 78:22]
  wire  bore_ldReq_0; // @[memGenTopLevel.scala 78:22]
  wire  bore_hitLD_0; // @[memGenTopLevel.scala 78:22]
  wire  bore_missLD_0; // @[memGenTopLevel.scala 78:22]
  wire  bore_cpuReq_0; // @[memGenTopLevel.scala 78:22]
  memoryWrapper memCtrl ( // @[memGenTopLevel.scala 67:25]
    .clock(memCtrl_clock),
    .reset(memCtrl_reset),
    .io_in_ready(memCtrl_io_in_ready),
    .io_in_valid(memCtrl_io_in_valid),
    .io_in_bits_addr(memCtrl_io_in_bits_addr),
    .io_in_bits_inst(memCtrl_io_in_bits_inst),
    .io_in_bits_data(memCtrl_io_in_bits_data),
    .io_in_bits_src(memCtrl_io_in_bits_src),
    .io_mem_aw_ready(memCtrl_io_mem_aw_ready),
    .io_mem_aw_valid(memCtrl_io_mem_aw_valid),
    .io_mem_aw_bits_addr(memCtrl_io_mem_aw_bits_addr),
    .io_mem_w_ready(memCtrl_io_mem_w_ready),
    .io_mem_w_valid(memCtrl_io_mem_w_valid),
    .io_mem_w_bits_data(memCtrl_io_mem_w_bits_data),
    .io_mem_b_ready(memCtrl_io_mem_b_ready),
    .io_mem_ar_ready(memCtrl_io_mem_ar_ready),
    .io_mem_ar_valid(memCtrl_io_mem_ar_valid),
    .io_mem_ar_bits_addr(memCtrl_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(memCtrl_io_mem_ar_bits_len),
    .io_mem_r_ready(memCtrl_io_mem_r_ready),
    .io_mem_r_valid(memCtrl_io_mem_r_valid),
    .io_mem_r_bits_data(memCtrl_io_mem_r_bits_data),
    .io_mem_r_bits_last(memCtrl_io_mem_r_bits_last),
    .io_out_ready(memCtrl_io_out_ready),
    .io_out_valid(memCtrl_io_out_valid),
    .io_out_bits_addr(memCtrl_io_out_bits_addr),
    .io_out_bits_data(memCtrl_io_out_bits_data),
    .io_out_bits_dst(memCtrl_io_out_bits_dst)
  );
  Queue memCtrlInputQueue ( // @[memGenTopLevel.scala 68:35]
    .clock(memCtrlInputQueue_clock),
    .reset(memCtrlInputQueue_reset),
    .io_enq_ready(memCtrlInputQueue_io_enq_ready),
    .io_enq_valid(memCtrlInputQueue_io_enq_valid),
    .io_enq_bits_addr(memCtrlInputQueue_io_enq_bits_addr),
    .io_enq_bits_inst(memCtrlInputQueue_io_enq_bits_inst),
    .io_enq_bits_data(memCtrlInputQueue_io_enq_bits_data),
    .io_enq_bits_src(memCtrlInputQueue_io_enq_bits_src),
    .io_deq_ready(memCtrlInputQueue_io_deq_ready),
    .io_deq_valid(memCtrlInputQueue_io_deq_valid),
    .io_deq_bits_addr(memCtrlInputQueue_io_deq_bits_addr),
    .io_deq_bits_inst(memCtrlInputQueue_io_deq_bits_inst),
    .io_deq_bits_data(memCtrlInputQueue_io_deq_bits_data),
    .io_deq_bits_src(memCtrlInputQueue_io_deq_bits_src)
  );
  Router routerNode_0 ( // @[memGenTopLevel.scala 70:28]
    .clock(routerNode_0_clock),
    .reset(routerNode_0_reset),
    .io_cacheIn_valid(routerNode_0_io_cacheIn_valid),
    .io_cacheIn_bits_addr(routerNode_0_io_cacheIn_bits_addr),
    .io_cacheIn_bits_inst(routerNode_0_io_cacheIn_bits_inst),
    .io_cacheIn_bits_data(routerNode_0_io_cacheIn_bits_data),
    .io_cacheOut_ready(routerNode_0_io_cacheOut_ready),
    .io_cacheOut_valid(routerNode_0_io_cacheOut_valid),
    .io_cacheOut_bits_addr(routerNode_0_io_cacheOut_bits_addr),
    .io_cacheOut_bits_inst(routerNode_0_io_cacheOut_bits_inst),
    .io_cacheOut_bits_data(routerNode_0_io_cacheOut_bits_data),
    .io_cacheOut_bits_msgType(routerNode_0_io_cacheOut_bits_msgType),
    .io_in_ready(routerNode_0_io_in_ready),
    .io_in_valid(routerNode_0_io_in_valid),
    .io_in_bits_addr(routerNode_0_io_in_bits_addr),
    .io_in_bits_inst(routerNode_0_io_in_bits_inst),
    .io_in_bits_data(routerNode_0_io_in_bits_data),
    .io_in_bits_src(routerNode_0_io_in_bits_src),
    .io_in_bits_dst(routerNode_0_io_in_bits_dst),
    .io_in_bits_msgType(routerNode_0_io_in_bits_msgType),
    .io_out_ready(routerNode_0_io_out_ready),
    .io_out_valid(routerNode_0_io_out_valid),
    .io_out_bits_addr(routerNode_0_io_out_bits_addr),
    .io_out_bits_inst(routerNode_0_io_out_bits_inst),
    .io_out_bits_data(routerNode_0_io_out_bits_data),
    .io_out_bits_src(routerNode_0_io_out_bits_src),
    .io_out_bits_dst(routerNode_0_io_out_bits_dst),
    .io_out_bits_msgType(routerNode_0_io_out_bits_msgType)
  );
  Router_1 routerNode_1 ( // @[memGenTopLevel.scala 70:28]
    .clock(routerNode_1_clock),
    .reset(routerNode_1_reset),
    .io_cacheIn_ready(routerNode_1_io_cacheIn_ready),
    .io_cacheIn_valid(routerNode_1_io_cacheIn_valid),
    .io_cacheIn_bits_addr(routerNode_1_io_cacheIn_bits_addr),
    .io_cacheIn_bits_data(routerNode_1_io_cacheIn_bits_data),
    .io_cacheIn_bits_dst(routerNode_1_io_cacheIn_bits_dst),
    .io_cacheOut_ready(routerNode_1_io_cacheOut_ready),
    .io_cacheOut_valid(routerNode_1_io_cacheOut_valid),
    .io_cacheOut_bits_addr(routerNode_1_io_cacheOut_bits_addr),
    .io_cacheOut_bits_inst(routerNode_1_io_cacheOut_bits_inst),
    .io_cacheOut_bits_data(routerNode_1_io_cacheOut_bits_data),
    .io_cacheOut_bits_src(routerNode_1_io_cacheOut_bits_src),
    .io_in_ready(routerNode_1_io_in_ready),
    .io_in_valid(routerNode_1_io_in_valid),
    .io_in_bits_addr(routerNode_1_io_in_bits_addr),
    .io_in_bits_inst(routerNode_1_io_in_bits_inst),
    .io_in_bits_data(routerNode_1_io_in_bits_data),
    .io_in_bits_src(routerNode_1_io_in_bits_src),
    .io_in_bits_dst(routerNode_1_io_in_bits_dst),
    .io_in_bits_msgType(routerNode_1_io_in_bits_msgType),
    .io_out_ready(routerNode_1_io_out_ready),
    .io_out_valid(routerNode_1_io_out_valid),
    .io_out_bits_addr(routerNode_1_io_out_bits_addr),
    .io_out_bits_inst(routerNode_1_io_out_bits_inst),
    .io_out_bits_data(routerNode_1_io_out_bits_data),
    .io_out_bits_src(routerNode_1_io_out_bits_src),
    .io_out_bits_dst(routerNode_1_io_out_bits_dst),
    .io_out_bits_msgType(routerNode_1_io_out_bits_msgType)
  );
  CacheNode cacheNode_0 ( // @[memGenTopLevel.scala 74:28]
    .clock(cacheNode_0_clock),
    .reset(cacheNode_0_reset),
    .io_in_cpu_ready(cacheNode_0_io_in_cpu_ready),
    .io_in_cpu_valid(cacheNode_0_io_in_cpu_valid),
    .io_in_cpu_bits_addr(cacheNode_0_io_in_cpu_bits_addr),
    .io_in_cpu_bits_inst(cacheNode_0_io_in_cpu_bits_inst),
    .io_in_cpu_bits_data(cacheNode_0_io_in_cpu_bits_data),
    .io_in_network_ready(cacheNode_0_io_in_network_ready),
    .io_in_network_valid(cacheNode_0_io_in_network_valid),
    .io_in_network_bits_addr(cacheNode_0_io_in_network_bits_addr),
    .io_in_network_bits_inst(cacheNode_0_io_in_network_bits_inst),
    .io_in_network_bits_data(cacheNode_0_io_in_network_bits_data),
    .io_in_network_bits_msgType(cacheNode_0_io_in_network_bits_msgType),
    .io_out_network_valid(cacheNode_0_io_out_network_valid),
    .io_out_network_bits_addr(cacheNode_0_io_out_network_bits_addr),
    .io_out_network_bits_inst(cacheNode_0_io_out_network_bits_inst),
    .io_out_network_bits_data(cacheNode_0_io_out_network_bits_data),
    .io_out_cpu_valid(cacheNode_0_io_out_cpu_valid),
    .io_out_cpu_bits_addr(cacheNode_0_io_out_cpu_bits_addr),
    ._T_814(cacheNode_0__T_814),
    ._T_808(cacheNode_0__T_808),
    ._T_819(cacheNode_0__T_819),
    .hitLD(cacheNode_0_hitLD),
    .missLD(cacheNode_0_missLD),
    ._T_811(cacheNode_0__T_811)
  );
  Bore bore ( // @[memGenTopLevel.scala 78:22]
    .clock(bore_clock),
    .reset(bore_reset),
    .io_events_0(bore_io_events_0),
    .io_events_1(bore_io_events_1),
    .io_events_2(bore_io_events_2),
    .io_events_3(bore_io_events_3),
    .io_events_4(bore_io_events_4),
    .io_events_5(bore_io_events_5),
    .memCtrlReq_0(bore_memCtrlReq_0),
    .instCount_0(bore_instCount_0),
    .ldReq_0(bore_ldReq_0),
    .hitLD_0(bore_hitLD_0),
    .missLD_0(bore_missLD_0),
    .cpuReq_0(bore_cpuReq_0)
  );
  assign io_instruction_0_ready = cacheNode_0_io_in_cpu_ready; // @[memGenTopLevel.scala 88:33]
  assign io_resp_0_valid = cacheNode_0_io_out_cpu_valid; // @[memGenTopLevel.scala 89:20]
  assign io_resp_0_bits_addr = cacheNode_0_io_out_cpu_bits_addr; // @[memGenTopLevel.scala 89:20]
  assign io_events_bits_0 = bore_io_events_0; // @[memGenTopLevel.scala 82:20]
  assign io_events_bits_1 = bore_io_events_1; // @[memGenTopLevel.scala 82:20]
  assign io_events_bits_2 = bore_io_events_2; // @[memGenTopLevel.scala 82:20]
  assign io_events_bits_3 = bore_io_events_3; // @[memGenTopLevel.scala 82:20]
  assign io_events_bits_4 = bore_io_events_4; // @[memGenTopLevel.scala 82:20]
  assign io_events_bits_5 = bore_io_events_5; // @[memGenTopLevel.scala 82:20]
  assign io_mem_aw_valid = memCtrl_io_mem_aw_valid; // @[memGenTopLevel.scala 100:12]
  assign io_mem_aw_bits_addr = memCtrl_io_mem_aw_bits_addr; // @[memGenTopLevel.scala 100:12]
  assign io_mem_w_valid = memCtrl_io_mem_w_valid; // @[memGenTopLevel.scala 100:12]
  assign io_mem_w_bits_data = memCtrl_io_mem_w_bits_data; // @[memGenTopLevel.scala 100:12]
  assign io_mem_b_ready = memCtrl_io_mem_b_ready; // @[memGenTopLevel.scala 100:12]
  assign io_mem_ar_valid = memCtrl_io_mem_ar_valid; // @[memGenTopLevel.scala 100:12]
  assign io_mem_ar_bits_addr = memCtrl_io_mem_ar_bits_addr; // @[memGenTopLevel.scala 100:12]
  assign io_mem_ar_bits_len = memCtrl_io_mem_ar_bits_len; // @[memGenTopLevel.scala 100:12]
  assign io_mem_r_ready = memCtrl_io_mem_r_ready; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_clock = clock;
  assign memCtrl_reset = reset;
  assign memCtrl_io_in_valid = memCtrlInputQueue_io_deq_valid; // @[memGenTopLevel.scala 98:19]
  assign memCtrl_io_in_bits_addr = memCtrlInputQueue_io_deq_bits_addr; // @[memGenTopLevel.scala 98:19]
  assign memCtrl_io_in_bits_inst = memCtrlInputQueue_io_deq_bits_inst; // @[memGenTopLevel.scala 98:19]
  assign memCtrl_io_in_bits_data = memCtrlInputQueue_io_deq_bits_data; // @[memGenTopLevel.scala 98:19]
  assign memCtrl_io_in_bits_src = memCtrlInputQueue_io_deq_bits_src; // @[memGenTopLevel.scala 98:19]
  assign memCtrl_io_mem_aw_ready = io_mem_aw_ready; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_io_mem_w_ready = io_mem_w_ready; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_io_mem_ar_ready = io_mem_ar_ready; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_io_mem_r_valid = io_mem_r_valid; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_io_mem_r_bits_data = io_mem_r_bits_data; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_io_mem_r_bits_last = io_mem_r_bits_last; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_io_out_ready = routerNode_1_io_cacheIn_ready; // @[memGenTopLevel.scala 99:52]
  assign memCtrlInputQueue_clock = clock;
  assign memCtrlInputQueue_reset = reset;
  assign memCtrlInputQueue_io_enq_valid = routerNode_1_io_cacheOut_valid; // @[memGenTopLevel.scala 97:30]
  assign memCtrlInputQueue_io_enq_bits_addr = routerNode_1_io_cacheOut_bits_addr; // @[memGenTopLevel.scala 97:30]
  assign memCtrlInputQueue_io_enq_bits_inst = routerNode_1_io_cacheOut_bits_inst; // @[memGenTopLevel.scala 97:30]
  assign memCtrlInputQueue_io_enq_bits_data = routerNode_1_io_cacheOut_bits_data; // @[memGenTopLevel.scala 97:30]
  assign memCtrlInputQueue_io_enq_bits_src = routerNode_1_io_cacheOut_bits_src; // @[memGenTopLevel.scala 97:30]
  assign memCtrlInputQueue_io_deq_ready = memCtrl_io_in_ready; // @[memGenTopLevel.scala 98:19]
  assign routerNode_0_clock = clock;
  assign routerNode_0_reset = reset;
  assign routerNode_0_io_cacheIn_valid = cacheNode_0_io_out_network_valid; // @[memGenTopLevel.scala 93:34]
  assign routerNode_0_io_cacheIn_bits_addr = cacheNode_0_io_out_network_bits_addr; // @[memGenTopLevel.scala 93:34]
  assign routerNode_0_io_cacheIn_bits_inst = cacheNode_0_io_out_network_bits_inst; // @[memGenTopLevel.scala 93:34]
  assign routerNode_0_io_cacheIn_bits_data = cacheNode_0_io_out_network_bits_data; // @[memGenTopLevel.scala 93:34]
  assign routerNode_0_io_cacheOut_ready = cacheNode_0_io_in_network_ready; // @[memGenTopLevel.scala 94:36]
  assign routerNode_0_io_in_valid = routerNode_1_io_out_valid; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_in_bits_addr = routerNode_1_io_out_bits_addr; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_in_bits_inst = routerNode_1_io_out_bits_inst; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_in_bits_data = routerNode_1_io_out_bits_data; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_in_bits_src = routerNode_1_io_out_bits_src; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_in_bits_dst = routerNode_1_io_out_bits_dst; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_in_bits_msgType = routerNode_1_io_out_bits_msgType; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_out_ready = routerNode_1_io_in_ready; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_clock = clock;
  assign routerNode_1_reset = reset;
  assign routerNode_1_io_cacheIn_valid = memCtrl_io_out_valid; // @[memGenTopLevel.scala 99:52]
  assign routerNode_1_io_cacheIn_bits_addr = memCtrl_io_out_bits_addr; // @[memGenTopLevel.scala 99:52]
  assign routerNode_1_io_cacheIn_bits_data = memCtrl_io_out_bits_data; // @[memGenTopLevel.scala 99:52]
  assign routerNode_1_io_cacheIn_bits_dst = memCtrl_io_out_bits_dst; // @[memGenTopLevel.scala 99:52]
  assign routerNode_1_io_cacheOut_ready = memCtrlInputQueue_io_enq_ready; // @[memGenTopLevel.scala 97:30]
  assign routerNode_1_io_in_valid = routerNode_0_io_out_valid; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_in_bits_addr = routerNode_0_io_out_bits_addr; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_in_bits_inst = routerNode_0_io_out_bits_inst; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_in_bits_data = routerNode_0_io_out_bits_data; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_in_bits_src = routerNode_0_io_out_bits_src; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_in_bits_dst = routerNode_0_io_out_bits_dst; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_in_bits_msgType = routerNode_0_io_out_bits_msgType; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_out_ready = routerNode_0_io_in_ready; // @[memGenTopLevel.scala 105:25]
  assign cacheNode_0_clock = clock;
  assign cacheNode_0_reset = reset;
  assign cacheNode_0_io_in_cpu_valid = io_instruction_0_valid; // @[memGenTopLevel.scala 87:38]
  assign cacheNode_0_io_in_cpu_bits_addr = io_instruction_0_bits_addr; // @[memGenTopLevel.scala 86:34]
  assign cacheNode_0_io_in_cpu_bits_inst = io_instruction_0_bits_inst; // @[memGenTopLevel.scala 86:34]
  assign cacheNode_0_io_in_cpu_bits_data = io_instruction_0_bits_data; // @[memGenTopLevel.scala 86:34]
  assign cacheNode_0_io_in_network_valid = routerNode_0_io_cacheOut_valid; // @[memGenTopLevel.scala 94:36]
  assign cacheNode_0_io_in_network_bits_addr = routerNode_0_io_cacheOut_bits_addr; // @[memGenTopLevel.scala 94:36]
  assign cacheNode_0_io_in_network_bits_inst = routerNode_0_io_cacheOut_bits_inst; // @[memGenTopLevel.scala 94:36]
  assign cacheNode_0_io_in_network_bits_data = routerNode_0_io_cacheOut_bits_data; // @[memGenTopLevel.scala 94:36]
  assign cacheNode_0_io_in_network_bits_msgType = routerNode_0_io_cacheOut_bits_msgType; // @[memGenTopLevel.scala 94:36]
  assign bore_clock = clock;
  assign bore_reset = reset;
  assign bore_memCtrlReq_0 = cacheNode_0__T_814;
  assign bore_instCount_0 = cacheNode_0__T_808;
  assign bore_ldReq_0 = cacheNode_0__T_819;
  assign bore_hitLD_0 = cacheNode_0_hitLD;
  assign bore_missLD_0 = cacheNode_0_missLD;
  assign bore_cpuReq_0 = cacheNode_0__T_811;
endmodule
module Arbiter_6(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits = io_in_0_bits; // @[Arbiter.scala 124:15]
endmodule
module Queue_47(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram [0:15]; // @[Decoupled.scala 209:16]
  wire [31:0] ram__T_11_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram__T_11_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram__T_3_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram__T_3_en; // @[Decoupled.scala 209:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 29:33]
  reg [3:0] deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  _T_1 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _T_5 = enq_ptr_value + 4'h1; // @[Counter.scala 39:22]
  wire  _GEN_9 = io_deq_ready ? 1'h0 : _T_1; // @[Decoupled.scala 240:27]
  wire  do_enq = empty ? _GEN_9 : _T_1; // @[Decoupled.scala 237:18]
  wire [3:0] _T_7 = deq_ptr_value + 4'h1; // @[Counter.scala 39:22]
  wire  do_deq = empty ? 1'h0 : _T_2; // @[Decoupled.scala 237:18]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  wire  _T_9 = ~empty; // @[Decoupled.scala 231:19]
  wire  _T_10 = ~full; // @[Decoupled.scala 232:19]
  assign ram__T_11_addr = deq_ptr_value;
  assign ram__T_11_data = ram[ram__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram__T_3_data = io_enq_bits;
  assign ram__T_3_addr = enq_ptr_value;
  assign ram__T_3_mask = 1'h1;
  assign ram__T_3_en = empty ? _GEN_9 : _T_1;
  assign io_enq_ready = io_deq_ready | _T_10; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = io_enq_valid | _T_9; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits = empty ? io_enq_bits : ram__T_11_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_3_en & ram__T_3_mask) begin
      ram[ram__T_3_addr] <= ram__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 4'h0;
    end else if (do_enq) begin
      enq_ptr_value <= _T_5;
    end
    if (reset) begin
      deq_ptr_value <= 4'h0;
    end else if (do_deq) begin
      deq_ptr_value <= _T_7;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _T_1;
        end
      end else begin
        maybe_full <= _T_1;
      end
    end
  end
endmodule
module memGenAccel(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_dataVals_field2_data,
  input  [63:0] io_in_bits_dataVals_field1_data,
  input  [63:0] io_in_bits_dataVals_field0_data,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_data_field1_data,
  output [31:0] io_events_bits_0,
  output [31:0] io_events_bits_1,
  output [31:0] io_events_bits_2,
  output [31:0] io_events_bits_3,
  output [31:0] io_events_bits_4,
  output [31:0] io_events_bits_5,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output        io_mem_b_ready,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [15:0] io_mem_ar_bits_len,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last
);
  wire  accel_clock; // @[memGenCacheShell.scala 24:22]
  wire  accel_reset; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_instruction_0_ready; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_instruction_0_valid; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_instruction_0_bits_addr; // @[memGenCacheShell.scala 24:22]
  wire [7:0] accel_io_instruction_0_bits_inst; // @[memGenCacheShell.scala 24:22]
  wire [63:0] accel_io_instruction_0_bits_data; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_resp_0_valid; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_resp_0_bits_addr; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_events_bits_0; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_events_bits_1; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_events_bits_2; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_events_bits_3; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_events_bits_4; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_events_bits_5; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_aw_ready; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_aw_valid; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_mem_aw_bits_addr; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_w_ready; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_w_valid; // @[memGenCacheShell.scala 24:22]
  wire [63:0] accel_io_mem_w_bits_data; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_b_ready; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_ar_ready; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_ar_valid; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_mem_ar_bits_addr; // @[memGenCacheShell.scala 24:22]
  wire [15:0] accel_io_mem_ar_bits_len; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_r_ready; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_r_valid; // @[memGenCacheShell.scala 24:22]
  wire [63:0] accel_io_mem_r_bits_data; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_r_bits_last; // @[memGenCacheShell.scala 24:22]
  wire  outArb_io_in_0_ready; // @[memGenCacheShell.scala 33:22]
  wire  outArb_io_in_0_valid; // @[memGenCacheShell.scala 33:22]
  wire [31:0] outArb_io_in_0_bits; // @[memGenCacheShell.scala 33:22]
  wire  outArb_io_out_ready; // @[memGenCacheShell.scala 33:22]
  wire  outArb_io_out_valid; // @[memGenCacheShell.scala 33:22]
  wire [31:0] outArb_io_out_bits; // @[memGenCacheShell.scala 33:22]
  wire  outAddrQueue_0_clock; // @[memGenCacheShell.scala 36:19]
  wire  outAddrQueue_0_reset; // @[memGenCacheShell.scala 36:19]
  wire  outAddrQueue_0_io_enq_ready; // @[memGenCacheShell.scala 36:19]
  wire  outAddrQueue_0_io_enq_valid; // @[memGenCacheShell.scala 36:19]
  wire [31:0] outAddrQueue_0_io_enq_bits; // @[memGenCacheShell.scala 36:19]
  wire  outAddrQueue_0_io_deq_ready; // @[memGenCacheShell.scala 36:19]
  wire  outAddrQueue_0_io_deq_valid; // @[memGenCacheShell.scala 36:19]
  wire [31:0] outAddrQueue_0_io_deq_bits; // @[memGenCacheShell.scala 36:19]
  wire  _T = io_in_bits_dataVals_field0_data == 64'h4; // @[memGenCacheShell.scala 47:54]
  wire [63:0] _GEN_1 = _T ? 64'h0 : io_in_bits_dataVals_field0_data; // @[memGenCacheShell.scala 47:68]
  memGenTopLevel accel ( // @[memGenCacheShell.scala 24:22]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_instruction_0_ready(accel_io_instruction_0_ready),
    .io_instruction_0_valid(accel_io_instruction_0_valid),
    .io_instruction_0_bits_addr(accel_io_instruction_0_bits_addr),
    .io_instruction_0_bits_inst(accel_io_instruction_0_bits_inst),
    .io_instruction_0_bits_data(accel_io_instruction_0_bits_data),
    .io_resp_0_valid(accel_io_resp_0_valid),
    .io_resp_0_bits_addr(accel_io_resp_0_bits_addr),
    .io_events_bits_0(accel_io_events_bits_0),
    .io_events_bits_1(accel_io_events_bits_1),
    .io_events_bits_2(accel_io_events_bits_2),
    .io_events_bits_3(accel_io_events_bits_3),
    .io_events_bits_4(accel_io_events_bits_4),
    .io_events_bits_5(accel_io_events_bits_5),
    .io_mem_aw_ready(accel_io_mem_aw_ready),
    .io_mem_aw_valid(accel_io_mem_aw_valid),
    .io_mem_aw_bits_addr(accel_io_mem_aw_bits_addr),
    .io_mem_w_ready(accel_io_mem_w_ready),
    .io_mem_w_valid(accel_io_mem_w_valid),
    .io_mem_w_bits_data(accel_io_mem_w_bits_data),
    .io_mem_b_ready(accel_io_mem_b_ready),
    .io_mem_ar_ready(accel_io_mem_ar_ready),
    .io_mem_ar_valid(accel_io_mem_ar_valid),
    .io_mem_ar_bits_addr(accel_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(accel_io_mem_ar_bits_len),
    .io_mem_r_ready(accel_io_mem_r_ready),
    .io_mem_r_valid(accel_io_mem_r_valid),
    .io_mem_r_bits_data(accel_io_mem_r_bits_data),
    .io_mem_r_bits_last(accel_io_mem_r_bits_last)
  );
  Arbiter_6 outArb ( // @[memGenCacheShell.scala 33:22]
    .io_in_0_ready(outArb_io_in_0_ready),
    .io_in_0_valid(outArb_io_in_0_valid),
    .io_in_0_bits(outArb_io_in_0_bits),
    .io_out_ready(outArb_io_out_ready),
    .io_out_valid(outArb_io_out_valid),
    .io_out_bits(outArb_io_out_bits)
  );
  Queue_47 outAddrQueue_0 ( // @[memGenCacheShell.scala 36:19]
    .clock(outAddrQueue_0_clock),
    .reset(outAddrQueue_0_reset),
    .io_enq_ready(outAddrQueue_0_io_enq_ready),
    .io_enq_valid(outAddrQueue_0_io_enq_valid),
    .io_enq_bits(outAddrQueue_0_io_enq_bits),
    .io_deq_ready(outAddrQueue_0_io_deq_ready),
    .io_deq_valid(outAddrQueue_0_io_deq_valid),
    .io_deq_bits(outAddrQueue_0_io_deq_bits)
  );
  assign io_in_ready = accel_io_instruction_0_ready; // @[memGenCacheShell.scala 45:15 memGenCacheShell.scala 56:17]
  assign io_out_valid = outArb_io_out_valid; // @[memGenCacheShell.scala 74:16]
  assign io_out_bits_data_field1_data = outArb_io_out_bits; // @[memGenCacheShell.scala 75:35]
  assign io_events_bits_0 = accel_io_events_bits_0; // @[memGenCacheShell.scala 78:13]
  assign io_events_bits_1 = accel_io_events_bits_1; // @[memGenCacheShell.scala 78:13]
  assign io_events_bits_2 = accel_io_events_bits_2; // @[memGenCacheShell.scala 78:13]
  assign io_events_bits_3 = accel_io_events_bits_3; // @[memGenCacheShell.scala 78:13]
  assign io_events_bits_4 = accel_io_events_bits_4; // @[memGenCacheShell.scala 78:13]
  assign io_events_bits_5 = accel_io_events_bits_5; // @[memGenCacheShell.scala 78:13]
  assign io_mem_aw_valid = accel_io_mem_aw_valid; // @[memGenCacheShell.scala 80:10]
  assign io_mem_aw_bits_addr = accel_io_mem_aw_bits_addr; // @[memGenCacheShell.scala 80:10]
  assign io_mem_w_valid = accel_io_mem_w_valid; // @[memGenCacheShell.scala 80:10]
  assign io_mem_w_bits_data = accel_io_mem_w_bits_data; // @[memGenCacheShell.scala 80:10]
  assign io_mem_b_ready = accel_io_mem_b_ready; // @[memGenCacheShell.scala 80:10]
  assign io_mem_ar_valid = accel_io_mem_ar_valid; // @[memGenCacheShell.scala 80:10]
  assign io_mem_ar_bits_addr = accel_io_mem_ar_bits_addr; // @[memGenCacheShell.scala 80:10]
  assign io_mem_ar_bits_len = accel_io_mem_ar_bits_len; // @[memGenCacheShell.scala 80:10]
  assign io_mem_r_ready = accel_io_mem_r_ready; // @[memGenCacheShell.scala 80:10]
  assign accel_clock = clock;
  assign accel_reset = reset;
  assign accel_io_instruction_0_valid = io_in_valid; // @[memGenCacheShell.scala 39:41 memGenCacheShell.scala 57:41]
  assign accel_io_instruction_0_bits_addr = io_in_bits_dataVals_field1_data[31:0]; // @[memGenCacheShell.scala 41:45 memGenCacheShell.scala 58:45]
  assign accel_io_instruction_0_bits_inst = _GEN_1[7:0]; // @[memGenCacheShell.scala 40:45 memGenCacheShell.scala 50:47 memGenCacheShell.scala 52:49]
  assign accel_io_instruction_0_bits_data = io_in_bits_dataVals_field2_data; // @[memGenCacheShell.scala 42:45 memGenCacheShell.scala 59:45]
  assign accel_io_mem_aw_ready = io_mem_aw_ready; // @[memGenCacheShell.scala 80:10]
  assign accel_io_mem_w_ready = io_mem_w_ready; // @[memGenCacheShell.scala 80:10]
  assign accel_io_mem_ar_ready = io_mem_ar_ready; // @[memGenCacheShell.scala 80:10]
  assign accel_io_mem_r_valid = io_mem_r_valid; // @[memGenCacheShell.scala 80:10]
  assign accel_io_mem_r_bits_data = io_mem_r_bits_data; // @[memGenCacheShell.scala 80:10]
  assign accel_io_mem_r_bits_last = io_mem_r_bits_last; // @[memGenCacheShell.scala 80:10]
  assign outArb_io_in_0_valid = outAddrQueue_0_io_deq_valid; // @[memGenCacheShell.scala 71:21]
  assign outArb_io_in_0_bits = outAddrQueue_0_io_deq_bits; // @[memGenCacheShell.scala 71:21]
  assign outArb_io_out_ready = io_out_ready; // @[memGenCacheShell.scala 76:23]
  assign outAddrQueue_0_clock = clock;
  assign outAddrQueue_0_reset = reset;
  assign outAddrQueue_0_io_enq_valid = accel_io_resp_0_valid; // @[memGenCacheShell.scala 68:34]
  assign outAddrQueue_0_io_enq_bits = accel_io_resp_0_valid ? accel_io_resp_0_bits_addr : 32'h0; // @[memGenCacheShell.scala 67:33]
  assign outAddrQueue_0_io_deq_ready = outArb_io_in_0_ready; // @[memGenCacheShell.scala 71:21]
endmodule
module Queue_48(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_data
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_data [0:999999]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_11_data; // @[Decoupled.scala 209:16]
  wire [19:0] ram_data__T_11_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire [19:0] ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [19:0] enq_ptr_value; // @[Counter.scala 29:33]
  reg [19:0] deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  _T_1 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = enq_ptr_value == 20'hf423f; // @[Counter.scala 38:24]
  wire [19:0] _T_5 = enq_ptr_value + 20'h1; // @[Counter.scala 39:22]
  wire  _GEN_13 = io_deq_ready ? 1'h0 : _T_1; // @[Decoupled.scala 240:27]
  wire  do_enq = empty ? _GEN_13 : _T_1; // @[Decoupled.scala 237:18]
  wire  wrap_1 = deq_ptr_value == 20'hf423f; // @[Counter.scala 38:24]
  wire [19:0] _T_7 = deq_ptr_value + 20'h1; // @[Counter.scala 39:22]
  wire  do_deq = empty ? 1'h0 : _T_2; // @[Decoupled.scala 237:18]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  wire  _T_9 = ~empty; // @[Decoupled.scala 231:19]
  wire  _T_10 = ~full; // @[Decoupled.scala 232:19]
  assign ram_data__T_11_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_data__T_11_data = ram_data[ram_data__T_11_addr]; // @[Decoupled.scala 209:16]
  `else
  assign ram_data__T_11_data = ram_data__T_11_addr >= 20'hf4240 ? _RAND_1[63:0] : ram_data[ram_data__T_11_addr]; // @[Decoupled.scala 209:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = enq_ptr_value;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = empty ? _GEN_13 : _T_1;
  assign io_enq_ready = io_deq_ready | _T_10; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = io_enq_valid | _T_9; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data__T_11_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {2{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1000000; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 20'h0;
    end else if (do_enq) begin
      if (wrap) begin
        enq_ptr_value <= 20'h0;
      end else begin
        enq_ptr_value <= _T_5;
      end
    end
    if (reset) begin
      deq_ptr_value <= 20'h0;
    end else if (do_deq) begin
      if (wrap_1) begin
        deq_ptr_value <= 20'h0;
      end else begin
        deq_ptr_value <= _T_7;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _T_1;
        end
      end else begin
        maybe_full <= _T_1;
      end
    end
  end
endmodule
module memGenDCRCacheShell(
  input         clock,
  input         reset,
  output        io_host_aw_ready,
  input         io_host_aw_valid,
  input  [31:0] io_host_aw_bits_addr,
  output        io_host_w_ready,
  input         io_host_w_valid,
  input  [63:0] io_host_w_bits_data,
  input         io_host_b_ready,
  output        io_host_b_valid,
  output        io_host_ar_ready,
  input         io_host_ar_valid,
  input  [31:0] io_host_ar_bits_addr,
  input         io_host_r_ready,
  output        io_host_r_valid,
  output [63:0] io_host_r_bits_data,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  output [31:0] io_mem_aw_bits_len,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output        io_mem_w_bits_last,
  output        io_mem_b_ready,
  input         io_mem_b_valid,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [31:0] io_mem_ar_bits_len,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  vcr_clock; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_reset; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_aw_ready; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_aw_valid; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_host_aw_bits_addr; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_w_ready; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_w_valid; // @[memGenDCRCacheShell.scala 37:19]
  wire [63:0] vcr_io_host_w_bits_data; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_b_ready; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_b_valid; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_ar_ready; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_ar_valid; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_host_ar_bits_addr; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_r_ready; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_r_valid; // @[memGenDCRCacheShell.scala 37:19]
  wire [63:0] vcr_io_host_r_bits_data; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_dcr_launch; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_dcr_finish; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_dcr_ecnt_0_valid; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_0_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_1_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_2_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_3_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_4_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_5_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_6_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_vals_0; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ptrs_0; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ptrs_1; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ptrs_2; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ptrs_3; // @[memGenDCRCacheShell.scala 37:19]
  wire  dmem_clock; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_reset; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_aw_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_aw_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_w_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_w_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_w_bits_last; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_b_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_b_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_ar_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_ar_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [31:0] dmem_io_mem_ar_bits_addr; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_r_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_r_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [63:0] dmem_io_mem_r_bits_data; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_r_bits_last; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_0_cmd_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [31:0] dmem_io_dme_rd_0_cmd_bits_addr; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_0_data_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_0_data_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [63:0] dmem_io_dme_rd_0_data_bits; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_1_cmd_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [31:0] dmem_io_dme_rd_1_cmd_bits_addr; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_1_data_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_1_data_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [63:0] dmem_io_dme_rd_1_data_bits; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_2_cmd_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [31:0] dmem_io_dme_rd_2_cmd_bits_addr; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_2_data_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_2_data_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [63:0] dmem_io_dme_rd_2_data_bits; // @[memGenDCRCacheShell.scala 38:20]
  wire  accel_clock; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_reset; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_in_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_in_valid; // @[memGenDCRCacheShell.scala 40:21]
  wire [63:0] accel_io_in_bits_dataVals_field2_data; // @[memGenDCRCacheShell.scala 40:21]
  wire [63:0] accel_io_in_bits_dataVals_field1_data; // @[memGenDCRCacheShell.scala 40:21]
  wire [63:0] accel_io_in_bits_dataVals_field0_data; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_out_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_out_valid; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_out_bits_data_field1_data; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_events_bits_0; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_events_bits_1; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_events_bits_2; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_events_bits_3; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_events_bits_4; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_events_bits_5; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_aw_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_aw_valid; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_mem_aw_bits_addr; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_w_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_w_valid; // @[memGenDCRCacheShell.scala 40:21]
  wire [63:0] accel_io_mem_w_bits_data; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_b_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_ar_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_ar_valid; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_mem_ar_bits_addr; // @[memGenDCRCacheShell.scala 40:21]
  wire [15:0] accel_io_mem_ar_bits_len; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_r_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_r_valid; // @[memGenDCRCacheShell.scala 40:21]
  wire [63:0] accel_io_mem_r_bits_data; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_r_bits_last; // @[memGenDCRCacheShell.scala 40:21]
  wire  inputQ_0_clock; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_0_reset; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_0_io_enq_ready; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_0_io_enq_valid; // @[memGenDCRCacheShell.scala 113:25]
  wire [63:0] inputQ_0_io_enq_bits_data; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_0_io_deq_ready; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_0_io_deq_valid; // @[memGenDCRCacheShell.scala 113:25]
  wire [63:0] inputQ_0_io_deq_bits_data; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_1_clock; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_1_reset; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_1_io_enq_ready; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_1_io_enq_valid; // @[memGenDCRCacheShell.scala 113:25]
  wire [63:0] inputQ_1_io_enq_bits_data; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_1_io_deq_ready; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_1_io_deq_valid; // @[memGenDCRCacheShell.scala 113:25]
  wire [63:0] inputQ_1_io_deq_bits_data; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_2_clock; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_2_reset; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_2_io_enq_ready; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_2_io_enq_valid; // @[memGenDCRCacheShell.scala 113:25]
  wire [63:0] inputQ_2_io_enq_bits_data; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_2_io_deq_ready; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_2_io_deq_valid; // @[memGenDCRCacheShell.scala 113:25]
  wire [63:0] inputQ_2_io_deq_bits_data; // @[memGenDCRCacheShell.scala 113:25]
  reg [2:0] state; // @[memGenDCRCacheShell.scala 46:22]
  reg [31:0] cycles; // @[memGenDCRCacheShell.scala 47:23]
  wire  last = state == 3'h5; // @[memGenDCRCacheShell.scala 48:20]
  wire  is_busy = state == 3'h2; // @[memGenDCRCacheShell.scala 49:23]
  reg [31:0] lastCycle; // @[memGenDCRCacheShell.scala 53:21]
  reg [14:0] cycle; // @[Counter.scala 29:33]
  wire  _T_1 = cycle == 15'h752f; // @[Counter.scala 38:24]
  wire [14:0] _T_3 = cycle + 15'h1; // @[Counter.scala 39:22]
  wire  stopSim = last & _T_1; // @[Counter.scala 67:17]
  wire  _T_4 = state == 3'h0; // @[memGenDCRCacheShell.scala 74:128]
  reg [63:0] vals_0; // @[Reg.scala 27:20]
  reg [63:0] ptrs_0; // @[Reg.scala 27:20]
  wire  _T_76 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_77 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_78 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_79 = ~inputQ_0_io_deq_valid; // @[memGenDCRCacheShell.scala 173:37]
  wire  _T_80 = inputQ_0_io_deq_bits_data == 64'h2; // @[memGenDCRCacheShell.scala 175:54]
  wire  _T_83 = inputQ_0_io_deq_bits_data == 64'h4; // @[memGenDCRCacheShell.scala 178:53]
  wire  _T_84 = accel_io_in_ready & accel_io_in_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_27 = _T_83 | _T_84; // @[memGenDCRCacheShell.scala 178:66]
  wire  _GEN_30 = _T_80 ? 1'h0 : _GEN_27; // @[memGenDCRCacheShell.scala 175:68]
  wire  _GEN_33 = _T_79 ? 1'h0 : _GEN_30; // @[memGenDCRCacheShell.scala 173:93]
  wire  _T_87 = 3'h4 == state; // @[Conditional.scala 37:30]
  reg [19:0] ackCounter; // @[Counter.scala 29:33]
  wire [63:0] _GEN_111 = {{44'd0}, ackCounter}; // @[memGenDCRCacheShell.scala 190:26]
  wire  _T_88 = _GEN_111 >= inputQ_2_io_deq_bits_data; // @[memGenDCRCacheShell.scala 190:26]
  wire  _GEN_40 = _T_87 & _T_88; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_78 ? _GEN_33 : _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_46 = _T_77 ? 1'h0 : _GEN_42; // @[Conditional.scala 39:67]
  wire  _T_19 = ackCounter == 20'hf423f; // @[Counter.scala 38:24]
  wire [19:0] _T_21 = ackCounter + 20'h1; // @[Counter.scala 39:22]
  wire  _GEN_44 = _T_78 ? 1'h0 : _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_48 = _T_77 ? 1'h0 : _GEN_44; // @[Conditional.scala 39:67]
  wire  resetAckCounter = _T_76 ? 1'h0 : _GEN_48; // @[Conditional.scala 40:58]
  reg [31:0] fillCounter; // @[memGenDCRCacheShell.scala 79:28]
  wire  _T_22 = dmem_io_mem_r_ready & dmem_io_mem_r_valid; // @[Decoupled.scala 40:37]
  reg [31:0] _T_29; // @[memGenDCRCacheShell.scala 92:22]
  wire [63:0] _T_30 = vals_0 / 64'h1; // @[memGenDCRCacheShell.scala 92:50]
  wire [63:0] _T_32 = _T_30 - 64'h1; // @[memGenDCRCacheShell.scala 92:61]
  wire [63:0] _GEN_112 = {{32'd0}, _T_29}; // @[memGenDCRCacheShell.scala 92:36]
  wire  fillWrap = _GEN_112 == _T_32; // @[memGenDCRCacheShell.scala 92:36]
  wire  _T_23 = fillWrap & _T_22; // @[memGenDCRCacheShell.scala 85:18]
  wire  _T_24 = _T_23 & dmem_io_mem_r_bits_last; // @[memGenDCRCacheShell.scala 85:42]
  wire  _T_26 = _T_22 & dmem_io_mem_r_bits_last; // @[memGenDCRCacheShell.scala 87:35]
  wire [31:0] _T_28 = fillCounter + 32'h1; // @[memGenDCRCacheShell.scala 88:32]
  reg [1:0] numQ; // @[Counter.scala 29:33]
  wire [1:0] _T_40 = numQ + 2'h1; // @[Counter.scala 39:22]
  wire  _T_43 = numQ == 2'h2; // @[memGenDCRCacheShell.scala 95:72]
  wire  _T_44 = _T_26 & _T_43; // @[memGenDCRCacheShell.scala 95:64]
  wire  goToBusy = _T_44 & fillWrap; // @[memGenDCRCacheShell.scala 95:80]
  wire [31:0] _T_47 = cycles + 32'h1; // @[memGenDCRCacheShell.scala 100:22]
  wire  _T_48 = accel_io_out_ready & accel_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_50 = ~reset; // @[memGenDCRCacheShell.scala 107:13]
  wire [32:0] _T_53 = fillCounter * 32'h1; // @[memGenDCRCacheShell.scala 120:79]
  wire [36:0] _T_54 = _T_53 * 33'h8; // @[memGenDCRCacheShell.scala 120:89]
  wire [36:0] _GEN_113 = {{5'd0}, vcr_io_dcr_ptrs_1}; // @[memGenDCRCacheShell.scala 120:65]
  wire [36:0] _T_56 = _GEN_113 + _T_54; // @[memGenDCRCacheShell.scala 120:65]
  wire [36:0] _GEN_114 = {{5'd0}, vcr_io_dcr_ptrs_2}; // @[memGenDCRCacheShell.scala 120:65]
  wire [36:0] _T_61 = _GEN_114 + _T_54; // @[memGenDCRCacheShell.scala 120:65]
  wire [36:0] _GEN_115 = {{5'd0}, vcr_io_dcr_ptrs_3}; // @[memGenDCRCacheShell.scala 120:65]
  wire [36:0] _T_66 = _GEN_115 + _T_54; // @[memGenDCRCacheShell.scala 120:65]
  wire  _T_68 = state == 3'h1; // @[memGenDCRCacheShell.scala 131:47]
  wire  _GEN_116 = 2'h0 == numQ; // @[memGenDCRCacheShell.scala 131:36]
  wire  _GEN_117 = 2'h1 == numQ; // @[memGenDCRCacheShell.scala 131:36]
  wire  _GEN_118 = 2'h2 == numQ; // @[memGenDCRCacheShell.scala 131:36]
  wire  _T_73 = is_busy | last; // @[memGenDCRCacheShell.scala 155:33]
  wire  _T_74 = state == 3'h4; // @[memGenDCRCacheShell.scala 155:59]
  wire  _GEN_28 = _T_83 ? 1'h0 : 1'h1; // @[memGenDCRCacheShell.scala 178:66]
  wire  _GEN_31 = _T_80 ? 1'h0 : _GEN_28; // @[memGenDCRCacheShell.scala 175:68]
  wire  _GEN_34 = _T_79 ? 1'h0 : _GEN_31; // @[memGenDCRCacheShell.scala 173:93]
  wire  _T_89 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_43 = _T_78 & _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_47 = _T_77 ? 1'h0 : _GEN_43; // @[Conditional.scala 39:67]
  wire  _GEN_122 = ~_T_76; // @[memGenDCRCacheShell.scala 177:17]
  wire  _GEN_123 = ~_T_77; // @[memGenDCRCacheShell.scala 177:17]
  wire  _GEN_124 = _GEN_122 & _GEN_123; // @[memGenDCRCacheShell.scala 177:17]
  wire  _GEN_125 = _GEN_124 & _T_78; // @[memGenDCRCacheShell.scala 177:17]
  wire  _GEN_126 = ~_T_79; // @[memGenDCRCacheShell.scala 177:17]
  wire  _GEN_127 = _GEN_125 & _GEN_126; // @[memGenDCRCacheShell.scala 177:17]
  wire  _GEN_128 = _GEN_127 & _T_80; // @[memGenDCRCacheShell.scala 177:17]
  wire  _GEN_135 = ~_T_80; // @[memGenDCRCacheShell.scala 183:21]
  wire  _GEN_136 = _GEN_127 & _GEN_135; // @[memGenDCRCacheShell.scala 183:21]
  wire  _GEN_137 = ~_T_83; // @[memGenDCRCacheShell.scala 183:21]
  wire  _GEN_138 = _GEN_136 & _GEN_137; // @[memGenDCRCacheShell.scala 183:21]
  wire  _GEN_139 = _GEN_138 & _T_84; // @[memGenDCRCacheShell.scala 183:21]
  DCR vcr ( // @[memGenDCRCacheShell.scala 37:19]
    .clock(vcr_clock),
    .reset(vcr_reset),
    .io_host_aw_ready(vcr_io_host_aw_ready),
    .io_host_aw_valid(vcr_io_host_aw_valid),
    .io_host_aw_bits_addr(vcr_io_host_aw_bits_addr),
    .io_host_w_ready(vcr_io_host_w_ready),
    .io_host_w_valid(vcr_io_host_w_valid),
    .io_host_w_bits_data(vcr_io_host_w_bits_data),
    .io_host_b_ready(vcr_io_host_b_ready),
    .io_host_b_valid(vcr_io_host_b_valid),
    .io_host_ar_ready(vcr_io_host_ar_ready),
    .io_host_ar_valid(vcr_io_host_ar_valid),
    .io_host_ar_bits_addr(vcr_io_host_ar_bits_addr),
    .io_host_r_ready(vcr_io_host_r_ready),
    .io_host_r_valid(vcr_io_host_r_valid),
    .io_host_r_bits_data(vcr_io_host_r_bits_data),
    .io_dcr_launch(vcr_io_dcr_launch),
    .io_dcr_finish(vcr_io_dcr_finish),
    .io_dcr_ecnt_0_valid(vcr_io_dcr_ecnt_0_valid),
    .io_dcr_ecnt_0_bits(vcr_io_dcr_ecnt_0_bits),
    .io_dcr_ecnt_1_bits(vcr_io_dcr_ecnt_1_bits),
    .io_dcr_ecnt_2_bits(vcr_io_dcr_ecnt_2_bits),
    .io_dcr_ecnt_3_bits(vcr_io_dcr_ecnt_3_bits),
    .io_dcr_ecnt_4_bits(vcr_io_dcr_ecnt_4_bits),
    .io_dcr_ecnt_5_bits(vcr_io_dcr_ecnt_5_bits),
    .io_dcr_ecnt_6_bits(vcr_io_dcr_ecnt_6_bits),
    .io_dcr_vals_0(vcr_io_dcr_vals_0),
    .io_dcr_ptrs_0(vcr_io_dcr_ptrs_0),
    .io_dcr_ptrs_1(vcr_io_dcr_ptrs_1),
    .io_dcr_ptrs_2(vcr_io_dcr_ptrs_2),
    .io_dcr_ptrs_3(vcr_io_dcr_ptrs_3)
  );
  DME dmem ( // @[memGenDCRCacheShell.scala 38:20]
    .clock(dmem_clock),
    .reset(dmem_reset),
    .io_mem_aw_ready(dmem_io_mem_aw_ready),
    .io_mem_aw_valid(dmem_io_mem_aw_valid),
    .io_mem_w_ready(dmem_io_mem_w_ready),
    .io_mem_w_valid(dmem_io_mem_w_valid),
    .io_mem_w_bits_last(dmem_io_mem_w_bits_last),
    .io_mem_b_ready(dmem_io_mem_b_ready),
    .io_mem_b_valid(dmem_io_mem_b_valid),
    .io_mem_ar_ready(dmem_io_mem_ar_ready),
    .io_mem_ar_valid(dmem_io_mem_ar_valid),
    .io_mem_ar_bits_addr(dmem_io_mem_ar_bits_addr),
    .io_mem_r_ready(dmem_io_mem_r_ready),
    .io_mem_r_valid(dmem_io_mem_r_valid),
    .io_mem_r_bits_data(dmem_io_mem_r_bits_data),
    .io_mem_r_bits_last(dmem_io_mem_r_bits_last),
    .io_dme_rd_0_cmd_valid(dmem_io_dme_rd_0_cmd_valid),
    .io_dme_rd_0_cmd_bits_addr(dmem_io_dme_rd_0_cmd_bits_addr),
    .io_dme_rd_0_data_ready(dmem_io_dme_rd_0_data_ready),
    .io_dme_rd_0_data_valid(dmem_io_dme_rd_0_data_valid),
    .io_dme_rd_0_data_bits(dmem_io_dme_rd_0_data_bits),
    .io_dme_rd_1_cmd_valid(dmem_io_dme_rd_1_cmd_valid),
    .io_dme_rd_1_cmd_bits_addr(dmem_io_dme_rd_1_cmd_bits_addr),
    .io_dme_rd_1_data_ready(dmem_io_dme_rd_1_data_ready),
    .io_dme_rd_1_data_valid(dmem_io_dme_rd_1_data_valid),
    .io_dme_rd_1_data_bits(dmem_io_dme_rd_1_data_bits),
    .io_dme_rd_2_cmd_valid(dmem_io_dme_rd_2_cmd_valid),
    .io_dme_rd_2_cmd_bits_addr(dmem_io_dme_rd_2_cmd_bits_addr),
    .io_dme_rd_2_data_ready(dmem_io_dme_rd_2_data_ready),
    .io_dme_rd_2_data_valid(dmem_io_dme_rd_2_data_valid),
    .io_dme_rd_2_data_bits(dmem_io_dme_rd_2_data_bits)
  );
  memGenAccel accel ( // @[memGenDCRCacheShell.scala 40:21]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_in_ready(accel_io_in_ready),
    .io_in_valid(accel_io_in_valid),
    .io_in_bits_dataVals_field2_data(accel_io_in_bits_dataVals_field2_data),
    .io_in_bits_dataVals_field1_data(accel_io_in_bits_dataVals_field1_data),
    .io_in_bits_dataVals_field0_data(accel_io_in_bits_dataVals_field0_data),
    .io_out_ready(accel_io_out_ready),
    .io_out_valid(accel_io_out_valid),
    .io_out_bits_data_field1_data(accel_io_out_bits_data_field1_data),
    .io_events_bits_0(accel_io_events_bits_0),
    .io_events_bits_1(accel_io_events_bits_1),
    .io_events_bits_2(accel_io_events_bits_2),
    .io_events_bits_3(accel_io_events_bits_3),
    .io_events_bits_4(accel_io_events_bits_4),
    .io_events_bits_5(accel_io_events_bits_5),
    .io_mem_aw_ready(accel_io_mem_aw_ready),
    .io_mem_aw_valid(accel_io_mem_aw_valid),
    .io_mem_aw_bits_addr(accel_io_mem_aw_bits_addr),
    .io_mem_w_ready(accel_io_mem_w_ready),
    .io_mem_w_valid(accel_io_mem_w_valid),
    .io_mem_w_bits_data(accel_io_mem_w_bits_data),
    .io_mem_b_ready(accel_io_mem_b_ready),
    .io_mem_ar_ready(accel_io_mem_ar_ready),
    .io_mem_ar_valid(accel_io_mem_ar_valid),
    .io_mem_ar_bits_addr(accel_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(accel_io_mem_ar_bits_len),
    .io_mem_r_ready(accel_io_mem_r_ready),
    .io_mem_r_valid(accel_io_mem_r_valid),
    .io_mem_r_bits_data(accel_io_mem_r_bits_data),
    .io_mem_r_bits_last(accel_io_mem_r_bits_last)
  );
  Queue_48 inputQ_0 ( // @[memGenDCRCacheShell.scala 113:25]
    .clock(inputQ_0_clock),
    .reset(inputQ_0_reset),
    .io_enq_ready(inputQ_0_io_enq_ready),
    .io_enq_valid(inputQ_0_io_enq_valid),
    .io_enq_bits_data(inputQ_0_io_enq_bits_data),
    .io_deq_ready(inputQ_0_io_deq_ready),
    .io_deq_valid(inputQ_0_io_deq_valid),
    .io_deq_bits_data(inputQ_0_io_deq_bits_data)
  );
  Queue_48 inputQ_1 ( // @[memGenDCRCacheShell.scala 113:25]
    .clock(inputQ_1_clock),
    .reset(inputQ_1_reset),
    .io_enq_ready(inputQ_1_io_enq_ready),
    .io_enq_valid(inputQ_1_io_enq_valid),
    .io_enq_bits_data(inputQ_1_io_enq_bits_data),
    .io_deq_ready(inputQ_1_io_deq_ready),
    .io_deq_valid(inputQ_1_io_deq_valid),
    .io_deq_bits_data(inputQ_1_io_deq_bits_data)
  );
  Queue_48 inputQ_2 ( // @[memGenDCRCacheShell.scala 113:25]
    .clock(inputQ_2_clock),
    .reset(inputQ_2_reset),
    .io_enq_ready(inputQ_2_io_enq_ready),
    .io_enq_valid(inputQ_2_io_enq_valid),
    .io_enq_bits_data(inputQ_2_io_enq_bits_data),
    .io_deq_ready(inputQ_2_io_deq_ready),
    .io_deq_valid(inputQ_2_io_deq_valid),
    .io_deq_bits_data(inputQ_2_io_deq_bits_data)
  );
  assign io_host_aw_ready = vcr_io_host_aw_ready; // @[memGenDCRCacheShell.scala 214:11]
  assign io_host_w_ready = vcr_io_host_w_ready; // @[memGenDCRCacheShell.scala 214:11]
  assign io_host_b_valid = vcr_io_host_b_valid; // @[memGenDCRCacheShell.scala 214:11]
  assign io_host_ar_ready = vcr_io_host_ar_ready; // @[memGenDCRCacheShell.scala 214:11]
  assign io_host_r_valid = vcr_io_host_r_valid; // @[memGenDCRCacheShell.scala 214:11]
  assign io_host_r_bits_data = vcr_io_host_r_bits_data; // @[memGenDCRCacheShell.scala 214:11]
  assign io_mem_aw_valid = _T_68 ? dmem_io_mem_aw_valid : accel_io_mem_aw_valid; // @[memGenDCRCacheShell.scala 207:12 memGenDCRCacheShell.scala 210:13]
  assign io_mem_aw_bits_addr = _T_68 ? 32'h0 : accel_io_mem_aw_bits_addr; // @[memGenDCRCacheShell.scala 207:12 memGenDCRCacheShell.scala 210:13]
  assign io_mem_aw_bits_len = _T_68 ? 32'h0 : 32'h1; // @[memGenDCRCacheShell.scala 207:12 memGenDCRCacheShell.scala 210:13]
  assign io_mem_w_valid = _T_68 ? 1'h0 : accel_io_mem_w_valid; // @[memGenDCRCacheShell.scala 207:12 memGenDCRCacheShell.scala 210:13]
  assign io_mem_w_bits_data = _T_68 ? 64'h0 : accel_io_mem_w_bits_data; // @[memGenDCRCacheShell.scala 207:12 memGenDCRCacheShell.scala 210:13]
  assign io_mem_w_bits_last = _T_68 & dmem_io_mem_w_bits_last; // @[memGenDCRCacheShell.scala 207:12 memGenDCRCacheShell.scala 210:13]
  assign io_mem_b_ready = _T_68 ? dmem_io_mem_b_ready : accel_io_mem_b_ready; // @[memGenDCRCacheShell.scala 207:12 memGenDCRCacheShell.scala 210:13]
  assign io_mem_ar_valid = _T_68 ? dmem_io_mem_ar_valid : accel_io_mem_ar_valid; // @[memGenDCRCacheShell.scala 207:12 memGenDCRCacheShell.scala 210:13]
  assign io_mem_ar_bits_addr = _T_68 ? dmem_io_mem_ar_bits_addr : accel_io_mem_ar_bits_addr; // @[memGenDCRCacheShell.scala 207:12 memGenDCRCacheShell.scala 210:13]
  assign io_mem_ar_bits_len = _T_68 ? 32'h0 : {{16'd0}, accel_io_mem_ar_bits_len}; // @[memGenDCRCacheShell.scala 207:12 memGenDCRCacheShell.scala 210:13]
  assign io_mem_r_ready = _T_68 ? dmem_io_mem_r_ready : accel_io_mem_r_ready; // @[memGenDCRCacheShell.scala 207:12 memGenDCRCacheShell.scala 210:13]
  assign vcr_clock = clock;
  assign vcr_reset = reset;
  assign vcr_io_host_aw_valid = io_host_aw_valid; // @[memGenDCRCacheShell.scala 214:11]
  assign vcr_io_host_aw_bits_addr = io_host_aw_bits_addr; // @[memGenDCRCacheShell.scala 214:11]
  assign vcr_io_host_w_valid = io_host_w_valid; // @[memGenDCRCacheShell.scala 214:11]
  assign vcr_io_host_w_bits_data = io_host_w_bits_data; // @[memGenDCRCacheShell.scala 214:11]
  assign vcr_io_host_b_ready = io_host_b_ready; // @[memGenDCRCacheShell.scala 214:11]
  assign vcr_io_host_ar_valid = io_host_ar_valid; // @[memGenDCRCacheShell.scala 214:11]
  assign vcr_io_host_ar_bits_addr = io_host_ar_bits_addr; // @[memGenDCRCacheShell.scala 214:11]
  assign vcr_io_host_r_ready = io_host_r_ready; // @[memGenDCRCacheShell.scala 214:11]
  assign vcr_io_dcr_finish = last & stopSim; // @[memGenDCRCacheShell.scala 204:21]
  assign vcr_io_dcr_ecnt_0_valid = state == 3'h5; // @[memGenDCRCacheShell.scala 103:27]
  assign vcr_io_dcr_ecnt_0_bits = lastCycle; // @[memGenDCRCacheShell.scala 104:26]
  assign vcr_io_dcr_ecnt_1_bits = accel_io_events_bits_0; // @[memGenDCRCacheShell.scala 63:31]
  assign vcr_io_dcr_ecnt_2_bits = accel_io_events_bits_1; // @[memGenDCRCacheShell.scala 63:31]
  assign vcr_io_dcr_ecnt_3_bits = accel_io_events_bits_2; // @[memGenDCRCacheShell.scala 63:31]
  assign vcr_io_dcr_ecnt_4_bits = accel_io_events_bits_3; // @[memGenDCRCacheShell.scala 63:31]
  assign vcr_io_dcr_ecnt_5_bits = accel_io_events_bits_4; // @[memGenDCRCacheShell.scala 63:31]
  assign vcr_io_dcr_ecnt_6_bits = accel_io_events_bits_5; // @[memGenDCRCacheShell.scala 63:31]
  assign dmem_clock = clock;
  assign dmem_reset = reset;
  assign dmem_io_mem_aw_ready = io_mem_aw_ready; // @[memGenDCRCacheShell.scala 207:12]
  assign dmem_io_mem_w_ready = io_mem_w_ready; // @[memGenDCRCacheShell.scala 207:12]
  assign dmem_io_mem_b_valid = io_mem_b_valid; // @[memGenDCRCacheShell.scala 207:12]
  assign dmem_io_mem_ar_ready = io_mem_ar_ready; // @[memGenDCRCacheShell.scala 207:12]
  assign dmem_io_mem_r_valid = io_mem_r_valid; // @[memGenDCRCacheShell.scala 207:12]
  assign dmem_io_mem_r_bits_data = io_mem_r_bits_data; // @[memGenDCRCacheShell.scala 207:12]
  assign dmem_io_mem_r_bits_last = io_mem_r_bits_last; // @[memGenDCRCacheShell.scala 207:12]
  assign dmem_io_dme_rd_0_cmd_valid = _GEN_116 & _T_68; // @[memGenDCRCacheShell.scala 122:39 memGenDCRCacheShell.scala 131:36]
  assign dmem_io_dme_rd_0_cmd_bits_addr = _T_56[31:0]; // @[memGenDCRCacheShell.scala 120:39]
  assign dmem_io_dme_rd_0_data_ready = inputQ_0_io_enq_ready; // @[memGenDCRCacheShell.scala 123:36]
  assign dmem_io_dme_rd_1_cmd_valid = _GEN_117 & _T_68; // @[memGenDCRCacheShell.scala 122:39 memGenDCRCacheShell.scala 131:36]
  assign dmem_io_dme_rd_1_cmd_bits_addr = _T_61[31:0]; // @[memGenDCRCacheShell.scala 120:39]
  assign dmem_io_dme_rd_1_data_ready = inputQ_1_io_enq_ready; // @[memGenDCRCacheShell.scala 123:36]
  assign dmem_io_dme_rd_2_cmd_valid = _GEN_118 & _T_68; // @[memGenDCRCacheShell.scala 122:39 memGenDCRCacheShell.scala 131:36]
  assign dmem_io_dme_rd_2_cmd_bits_addr = _T_66[31:0]; // @[memGenDCRCacheShell.scala 120:39]
  assign dmem_io_dme_rd_2_data_ready = inputQ_2_io_enq_ready; // @[memGenDCRCacheShell.scala 123:36]
  assign accel_clock = clock;
  assign accel_reset = reset;
  assign accel_io_in_valid = _T_76 ? 1'h0 : _GEN_47; // @[memGenDCRCacheShell.scala 154:21 memGenDCRCacheShell.scala 181:31]
  assign accel_io_in_bits_dataVals_field2_data = inputQ_2_io_deq_bits_data; // @[memGenDCRCacheShell.scala 143:49]
  assign accel_io_in_bits_dataVals_field1_data = inputQ_1_io_deq_bits_data + ptrs_0; // @[memGenDCRCacheShell.scala 141:50]
  assign accel_io_in_bits_dataVals_field0_data = inputQ_0_io_deq_bits_data; // @[memGenDCRCacheShell.scala 143:49]
  assign accel_io_out_ready = _T_73 | _T_74; // @[memGenDCRCacheShell.scala 155:22]
  assign accel_io_mem_aw_ready = io_mem_aw_ready; // @[memGenDCRCacheShell.scala 210:13]
  assign accel_io_mem_w_ready = io_mem_w_ready; // @[memGenDCRCacheShell.scala 210:13]
  assign accel_io_mem_ar_ready = io_mem_ar_ready; // @[memGenDCRCacheShell.scala 210:13]
  assign accel_io_mem_r_valid = io_mem_r_valid; // @[memGenDCRCacheShell.scala 210:13]
  assign accel_io_mem_r_bits_data = io_mem_r_bits_data; // @[memGenDCRCacheShell.scala 210:13]
  assign accel_io_mem_r_bits_last = io_mem_r_bits_last; // @[memGenDCRCacheShell.scala 210:13]
  assign inputQ_0_clock = clock;
  assign inputQ_0_reset = reset;
  assign inputQ_0_io_enq_valid = dmem_io_dme_rd_0_data_valid; // @[memGenDCRCacheShell.scala 126:30]
  assign inputQ_0_io_enq_bits_data = dmem_io_dme_rd_0_data_bits; // @[memGenDCRCacheShell.scala 125:29]
  assign inputQ_0_io_deq_ready = _T_76 ? 1'h0 : _GEN_46; // @[memGenDCRCacheShell.scala 127:30]
  assign inputQ_1_clock = clock;
  assign inputQ_1_reset = reset;
  assign inputQ_1_io_enq_valid = dmem_io_dme_rd_1_data_valid; // @[memGenDCRCacheShell.scala 126:30]
  assign inputQ_1_io_enq_bits_data = dmem_io_dme_rd_1_data_bits; // @[memGenDCRCacheShell.scala 125:29]
  assign inputQ_1_io_deq_ready = _T_76 ? 1'h0 : _GEN_46; // @[memGenDCRCacheShell.scala 127:30]
  assign inputQ_2_clock = clock;
  assign inputQ_2_reset = reset;
  assign inputQ_2_io_enq_valid = dmem_io_dme_rd_2_data_valid; // @[memGenDCRCacheShell.scala 126:30]
  assign inputQ_2_io_enq_bits_data = dmem_io_dme_rd_2_data_bits; // @[memGenDCRCacheShell.scala 125:29]
  assign inputQ_2_io_deq_ready = _T_76 ? 1'h0 : _GEN_46; // @[memGenDCRCacheShell.scala 127:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  cycles = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  lastCycle = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  cycle = _RAND_3[14:0];
  _RAND_4 = {2{`RANDOM}};
  vals_0 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ptrs_0 = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  ackCounter = _RAND_6[19:0];
  _RAND_7 = {1{`RANDOM}};
  fillCounter = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _T_29 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  numQ = _RAND_9[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else if (_T_76) begin
      if (vcr_io_dcr_launch) begin
        state <= 3'h1;
      end
    end else if (_T_77) begin
      if (goToBusy) begin
        state <= 3'h2;
      end
    end else if (_T_78) begin
      if (_T_79) begin
        state <= 3'h5;
      end else if (_T_80) begin
        state <= 3'h4;
      end
    end else if (_T_87) begin
      if (_T_88) begin
        state <= 3'h2;
      end
    end else if (_T_89) begin
      if (stopSim) begin
        state <= 3'h0;
      end
    end
    if (reset) begin
      cycles <= 32'h0;
    end else if (goToBusy) begin
      cycles <= 32'h0;
    end else begin
      cycles <= _T_47;
    end
    if (_T_48) begin
      lastCycle <= cycles;
    end
    if (reset) begin
      cycle <= 15'h0;
    end else if (last) begin
      if (_T_1) begin
        cycle <= 15'h0;
      end else begin
        cycle <= _T_3;
      end
    end
    if (reset) begin
      vals_0 <= 64'h0;
    end else if (_T_4) begin
      vals_0 <= {{32'd0}, vcr_io_dcr_vals_0};
    end
    if (reset) begin
      ptrs_0 <= 64'h0;
    end else if (_T_4) begin
      ptrs_0 <= {{32'd0}, vcr_io_dcr_ptrs_0};
    end
    if (reset) begin
      ackCounter <= 20'h0;
    end else if (resetAckCounter) begin
      ackCounter <= 20'h0;
    end else if (accel_io_out_valid) begin
      if (_T_19) begin
        ackCounter <= 20'h0;
      end else begin
        ackCounter <= _T_21;
      end
    end
    if (reset) begin
      fillCounter <= 32'h0;
    end else if (_T_24) begin
      fillCounter <= 32'h0;
    end else if (_T_26) begin
      fillCounter <= _T_28;
    end
    _T_29 <= fillCounter;
    if (reset) begin
      numQ <= 2'h0;
    end else if (_T_24) begin
      numQ <= _T_40;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_48 & _T_50) begin
          $fwrite(32'h80000002,"Data back for addr %d cycle %d \n",accel_io_out_bits_data_field1_data,cycles); // @[memGenDCRCacheShell.scala 107:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_48 & _T_50) begin
          $fwrite(32'h80000002,"ackCounter :%d\n",ackCounter); // @[memGenDCRCacheShell.scala 108:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_128 & _T_50) begin
          $fwrite(32'h80000002,"Ack \n"); // @[memGenDCRCacheShell.scala 177:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_139 & _T_50) begin
          $fwrite(32'h80000002,"\nInst : %d for addr %d with data %d cycle %d \n",accel_io_in_bits_dataVals_field0_data,accel_io_in_bits_dataVals_field1_data,accel_io_in_bits_dataVals_field2_data,cycles); // @[memGenDCRCacheShell.scala 183:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module DandelionSimDCRAccel(
  input   clock,
  input   reset,
  input   sim_clock,
  output  sim_wait
);
  wire  sim_shell_clock; // @[DCRAccel.scala 52:25]
  wire  sim_shell_reset; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_aw_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_aw_valid; // @[DCRAccel.scala 52:25]
  wire [31:0] sim_shell_mem_aw_bits_addr; // @[DCRAccel.scala 52:25]
  wire [31:0] sim_shell_mem_aw_bits_len; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_w_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_w_valid; // @[DCRAccel.scala 52:25]
  wire [63:0] sim_shell_mem_w_bits_data; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_w_bits_last; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_b_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_b_valid; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_ar_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_ar_valid; // @[DCRAccel.scala 52:25]
  wire [31:0] sim_shell_mem_ar_bits_addr; // @[DCRAccel.scala 52:25]
  wire [31:0] sim_shell_mem_ar_bits_len; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_r_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_r_valid; // @[DCRAccel.scala 52:25]
  wire [63:0] sim_shell_mem_r_bits_data; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_r_bits_last; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_aw_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_aw_valid; // @[DCRAccel.scala 52:25]
  wire [31:0] sim_shell_host_aw_bits_addr; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_w_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_w_valid; // @[DCRAccel.scala 52:25]
  wire [63:0] sim_shell_host_w_bits_data; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_b_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_b_valid; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_ar_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_ar_valid; // @[DCRAccel.scala 52:25]
  wire [31:0] sim_shell_host_ar_bits_addr; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_r_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_r_valid; // @[DCRAccel.scala 52:25]
  wire [63:0] sim_shell_host_r_bits_data; // @[DCRAccel.scala 52:25]
  wire  sim_shell_sim_clock; // @[DCRAccel.scala 52:25]
  wire  sim_shell_sim_wait; // @[DCRAccel.scala 52:25]
  wire  shell_clock; // @[DCRAccel.scala 53:21]
  wire  shell_reset; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_aw_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_aw_valid; // @[DCRAccel.scala 53:21]
  wire [31:0] shell_io_host_aw_bits_addr; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_w_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_w_valid; // @[DCRAccel.scala 53:21]
  wire [63:0] shell_io_host_w_bits_data; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_b_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_b_valid; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_ar_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_ar_valid; // @[DCRAccel.scala 53:21]
  wire [31:0] shell_io_host_ar_bits_addr; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_r_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_r_valid; // @[DCRAccel.scala 53:21]
  wire [63:0] shell_io_host_r_bits_data; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_aw_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_aw_valid; // @[DCRAccel.scala 53:21]
  wire [31:0] shell_io_mem_aw_bits_addr; // @[DCRAccel.scala 53:21]
  wire [31:0] shell_io_mem_aw_bits_len; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_w_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_w_valid; // @[DCRAccel.scala 53:21]
  wire [63:0] shell_io_mem_w_bits_data; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_w_bits_last; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_b_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_b_valid; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_ar_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_ar_valid; // @[DCRAccel.scala 53:21]
  wire [31:0] shell_io_mem_ar_bits_addr; // @[DCRAccel.scala 53:21]
  wire [31:0] shell_io_mem_ar_bits_len; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_r_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_r_valid; // @[DCRAccel.scala 53:21]
  wire [63:0] shell_io_mem_r_bits_data; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_r_bits_last; // @[DCRAccel.scala 53:21]
  AXISimShell sim_shell ( // @[DCRAccel.scala 52:25]
    .clock(sim_shell_clock),
    .reset(sim_shell_reset),
    .mem_aw_ready(sim_shell_mem_aw_ready),
    .mem_aw_valid(sim_shell_mem_aw_valid),
    .mem_aw_bits_addr(sim_shell_mem_aw_bits_addr),
    .mem_aw_bits_len(sim_shell_mem_aw_bits_len),
    .mem_w_ready(sim_shell_mem_w_ready),
    .mem_w_valid(sim_shell_mem_w_valid),
    .mem_w_bits_data(sim_shell_mem_w_bits_data),
    .mem_w_bits_last(sim_shell_mem_w_bits_last),
    .mem_b_ready(sim_shell_mem_b_ready),
    .mem_b_valid(sim_shell_mem_b_valid),
    .mem_ar_ready(sim_shell_mem_ar_ready),
    .mem_ar_valid(sim_shell_mem_ar_valid),
    .mem_ar_bits_addr(sim_shell_mem_ar_bits_addr),
    .mem_ar_bits_len(sim_shell_mem_ar_bits_len),
    .mem_r_ready(sim_shell_mem_r_ready),
    .mem_r_valid(sim_shell_mem_r_valid),
    .mem_r_bits_data(sim_shell_mem_r_bits_data),
    .mem_r_bits_last(sim_shell_mem_r_bits_last),
    .host_aw_ready(sim_shell_host_aw_ready),
    .host_aw_valid(sim_shell_host_aw_valid),
    .host_aw_bits_addr(sim_shell_host_aw_bits_addr),
    .host_w_ready(sim_shell_host_w_ready),
    .host_w_valid(sim_shell_host_w_valid),
    .host_w_bits_data(sim_shell_host_w_bits_data),
    .host_b_ready(sim_shell_host_b_ready),
    .host_b_valid(sim_shell_host_b_valid),
    .host_ar_ready(sim_shell_host_ar_ready),
    .host_ar_valid(sim_shell_host_ar_valid),
    .host_ar_bits_addr(sim_shell_host_ar_bits_addr),
    .host_r_ready(sim_shell_host_r_ready),
    .host_r_valid(sim_shell_host_r_valid),
    .host_r_bits_data(sim_shell_host_r_bits_data),
    .sim_clock(sim_shell_sim_clock),
    .sim_wait(sim_shell_sim_wait)
  );
  memGenDCRCacheShell shell ( // @[DCRAccel.scala 53:21]
    .clock(shell_clock),
    .reset(shell_reset),
    .io_host_aw_ready(shell_io_host_aw_ready),
    .io_host_aw_valid(shell_io_host_aw_valid),
    .io_host_aw_bits_addr(shell_io_host_aw_bits_addr),
    .io_host_w_ready(shell_io_host_w_ready),
    .io_host_w_valid(shell_io_host_w_valid),
    .io_host_w_bits_data(shell_io_host_w_bits_data),
    .io_host_b_ready(shell_io_host_b_ready),
    .io_host_b_valid(shell_io_host_b_valid),
    .io_host_ar_ready(shell_io_host_ar_ready),
    .io_host_ar_valid(shell_io_host_ar_valid),
    .io_host_ar_bits_addr(shell_io_host_ar_bits_addr),
    .io_host_r_ready(shell_io_host_r_ready),
    .io_host_r_valid(shell_io_host_r_valid),
    .io_host_r_bits_data(shell_io_host_r_bits_data),
    .io_mem_aw_ready(shell_io_mem_aw_ready),
    .io_mem_aw_valid(shell_io_mem_aw_valid),
    .io_mem_aw_bits_addr(shell_io_mem_aw_bits_addr),
    .io_mem_aw_bits_len(shell_io_mem_aw_bits_len),
    .io_mem_w_ready(shell_io_mem_w_ready),
    .io_mem_w_valid(shell_io_mem_w_valid),
    .io_mem_w_bits_data(shell_io_mem_w_bits_data),
    .io_mem_w_bits_last(shell_io_mem_w_bits_last),
    .io_mem_b_ready(shell_io_mem_b_ready),
    .io_mem_b_valid(shell_io_mem_b_valid),
    .io_mem_ar_ready(shell_io_mem_ar_ready),
    .io_mem_ar_valid(shell_io_mem_ar_valid),
    .io_mem_ar_bits_addr(shell_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(shell_io_mem_ar_bits_len),
    .io_mem_r_ready(shell_io_mem_r_ready),
    .io_mem_r_valid(shell_io_mem_r_valid),
    .io_mem_r_bits_data(shell_io_mem_r_bits_data),
    .io_mem_r_bits_last(shell_io_mem_r_bits_last)
  );
  assign sim_wait = sim_shell_sim_wait; // @[DCRAccel.scala 56:12]
  assign sim_shell_clock = clock;
  assign sim_shell_reset = reset;
  assign sim_shell_mem_aw_valid = shell_io_mem_aw_valid; // @[DCRAccel.scala 62:20]
  assign sim_shell_mem_aw_bits_addr = shell_io_mem_aw_bits_addr; // @[DCRAccel.scala 62:20]
  assign sim_shell_mem_aw_bits_len = shell_io_mem_aw_bits_len; // @[DCRAccel.scala 62:20]
  assign sim_shell_mem_w_valid = shell_io_mem_w_valid; // @[DCRAccel.scala 63:19]
  assign sim_shell_mem_w_bits_data = shell_io_mem_w_bits_data; // @[DCRAccel.scala 63:19]
  assign sim_shell_mem_w_bits_last = shell_io_mem_w_bits_last; // @[DCRAccel.scala 63:19]
  assign sim_shell_mem_b_ready = shell_io_mem_b_ready; // @[DCRAccel.scala 64:18]
  assign sim_shell_mem_ar_valid = shell_io_mem_ar_valid; // @[DCRAccel.scala 61:20]
  assign sim_shell_mem_ar_bits_addr = shell_io_mem_ar_bits_addr; // @[DCRAccel.scala 61:20]
  assign sim_shell_mem_ar_bits_len = shell_io_mem_ar_bits_len; // @[DCRAccel.scala 61:20]
  assign sim_shell_mem_r_ready = shell_io_mem_r_ready; // @[DCRAccel.scala 65:18]
  assign sim_shell_host_aw_ready = shell_io_host_aw_ready; // @[DCRAccel.scala 70:20]
  assign sim_shell_host_w_ready = shell_io_host_w_ready; // @[DCRAccel.scala 71:19]
  assign sim_shell_host_b_valid = shell_io_host_b_valid; // @[DCRAccel.scala 67:20]
  assign sim_shell_host_ar_ready = shell_io_host_ar_ready; // @[DCRAccel.scala 69:20]
  assign sim_shell_host_r_valid = shell_io_host_r_valid; // @[DCRAccel.scala 68:20]
  assign sim_shell_host_r_bits_data = shell_io_host_r_bits_data; // @[DCRAccel.scala 68:20]
  assign sim_shell_sim_clock = sim_clock; // @[DCRAccel.scala 55:23]
  assign shell_clock = clock;
  assign shell_reset = reset;
  assign shell_io_host_aw_valid = sim_shell_host_aw_valid; // @[DCRAccel.scala 70:20]
  assign shell_io_host_aw_bits_addr = sim_shell_host_aw_bits_addr; // @[DCRAccel.scala 70:20]
  assign shell_io_host_w_valid = sim_shell_host_w_valid; // @[DCRAccel.scala 71:19]
  assign shell_io_host_w_bits_data = sim_shell_host_w_bits_data; // @[DCRAccel.scala 71:19]
  assign shell_io_host_b_ready = sim_shell_host_b_ready; // @[DCRAccel.scala 67:20]
  assign shell_io_host_ar_valid = sim_shell_host_ar_valid; // @[DCRAccel.scala 69:20]
  assign shell_io_host_ar_bits_addr = sim_shell_host_ar_bits_addr; // @[DCRAccel.scala 69:20]
  assign shell_io_host_r_ready = sim_shell_host_r_ready; // @[DCRAccel.scala 68:20]
  assign shell_io_mem_aw_ready = sim_shell_mem_aw_ready; // @[DCRAccel.scala 62:20]
  assign shell_io_mem_w_ready = sim_shell_mem_w_ready; // @[DCRAccel.scala 63:19]
  assign shell_io_mem_b_valid = sim_shell_mem_b_valid; // @[DCRAccel.scala 64:18]
  assign shell_io_mem_ar_ready = sim_shell_mem_ar_ready; // @[DCRAccel.scala 61:20]
  assign shell_io_mem_r_valid = sim_shell_mem_r_valid; // @[DCRAccel.scala 65:18]
  assign shell_io_mem_r_bits_data = sim_shell_mem_r_bits_data; // @[DCRAccel.scala 65:18]
  assign shell_io_mem_r_bits_last = sim_shell_mem_r_bits_last; // @[DCRAccel.scala 65:18]
endmodule
