module VTASim(
  input   clock,
  input   reset,
  output  sim_wait
);
  wire  sim_clock; // @[SimShell.scala 55:19]
  wire  sim_reset; // @[SimShell.scala 55:19]
  wire  sim_dpi_wait; // @[SimShell.scala 55:19]
  VTASimDPI sim ( // @[SimShell.scala 55:19]
    .clock(sim_clock),
    .reset(sim_reset),
    .dpi_wait(sim_dpi_wait)
  );
  assign sim_wait = sim_dpi_wait; // @[SimShell.scala 58:12]
  assign sim_clock = clock; // @[SimShell.scala 57:16]
  assign sim_reset = reset; // @[SimShell.scala 56:16]
endmodule
module VTAHostDPIToAXI(
  input         clock,
  input         reset,
  input         io_dpi_req_valid,
  input         io_dpi_req_opcode,
  input  [31:0] io_dpi_req_addr,
  input  [31:0] io_dpi_req_value,
  output        io_dpi_req_deq,
  output        io_dpi_resp_valid,
  output [31:0] io_dpi_resp_bits,
  input         io_axi_aw_ready,
  output        io_axi_aw_valid,
  output [31:0] io_axi_aw_bits_addr,
  input         io_axi_w_ready,
  output        io_axi_w_valid,
  output [63:0] io_axi_w_bits_data,
  output        io_axi_b_ready,
  input         io_axi_b_valid,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [31:0] io_axi_ar_bits_addr,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [63:0] io_axi_r_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] addr; // @[VTAHostDPI.scala 69:21]
  reg [31:0] data; // @[VTAHostDPI.scala 70:21]
  reg [2:0] state; // @[VTAHostDPI.scala 73:22]
  wire  _T_2 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_6 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_8 = state == 3'h0; // @[VTAHostDPI.scala 112:14]
  wire  _T_9 = _T_8 & io_dpi_req_valid; // @[VTAHostDPI.scala 112:24]
  wire  _T_10 = state == 3'h3; // @[VTAHostDPI.scala 117:28]
  wire  _T_13 = state == 3'h1; // @[VTAHostDPI.scala 124:28]
  wire  _T_16 = _T_13 & io_axi_ar_ready; // @[VTAHostDPI.scala 128:45]
  wire  _T_18 = _T_10 & io_axi_aw_ready; // @[VTAHostDPI.scala 128:91]
  assign io_dpi_req_deq = _T_16 | _T_18; // @[VTAHostDPI.scala 128:18]
  assign io_dpi_resp_valid = io_axi_r_valid; // @[VTAHostDPI.scala 129:21]
  assign io_dpi_resp_bits = io_axi_r_bits_data[31:0]; // @[VTAHostDPI.scala 130:20]
  assign io_axi_aw_valid = state == 3'h3; // @[VTAHostDPI.scala 117:19]
  assign io_axi_aw_bits_addr = addr; // @[VTAHostDPI.scala 118:23]
  assign io_axi_w_valid = state == 3'h4; // @[VTAHostDPI.scala 119:18]
  assign io_axi_w_bits_data = {{32'd0}, data}; // @[VTAHostDPI.scala 120:22]
  assign io_axi_b_ready = state == 3'h5; // @[VTAHostDPI.scala 122:18]
  assign io_axi_ar_valid = state == 3'h1; // @[VTAHostDPI.scala 124:19]
  assign io_axi_ar_bits_addr = addr; // @[VTAHostDPI.scala 125:23]
  assign io_axi_r_ready = state == 3'h2; // @[VTAHostDPI.scala 126:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  data = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr <= 32'h0;
    end else if (_T_9) begin
      addr <= io_dpi_req_addr;
    end
    if (reset) begin
      data <= 32'h0;
    end else if (_T_9) begin
      data <= io_dpi_req_value;
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_2) begin
      if (io_dpi_req_valid) begin
        if (io_dpi_req_opcode) begin
          state <= 3'h3;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (_T_3) begin
      if (io_axi_ar_ready) begin
        state <= 3'h2;
      end
    end else if (_T_4) begin
      if (io_axi_r_valid) begin
        state <= 3'h0;
      end
    end else if (_T_5) begin
      if (io_axi_aw_ready) begin
        state <= 3'h4;
      end
    end else if (_T_6) begin
      if (io_axi_w_ready) begin
        state <= 3'h5;
      end
    end else if (_T_7) begin
      if (io_axi_b_valid) begin
        state <= 3'h0;
      end
    end
  end
endmodule
module VTAHost(
  input         clock,
  input         reset,
  input         io_axi_aw_ready,
  output        io_axi_aw_valid,
  output [31:0] io_axi_aw_bits_addr,
  input         io_axi_w_ready,
  output        io_axi_w_valid,
  output [63:0] io_axi_w_bits_data,
  output        io_axi_b_ready,
  input         io_axi_b_valid,
  input         io_axi_ar_ready,
  output        io_axi_ar_valid,
  output [31:0] io_axi_ar_bits_addr,
  output        io_axi_r_ready,
  input         io_axi_r_valid,
  input  [63:0] io_axi_r_bits_data
);
  wire  host_dpi_clock; // @[SimShell.scala 20:24]
  wire  host_dpi_reset; // @[SimShell.scala 20:24]
  wire  host_dpi_dpi_req_valid; // @[SimShell.scala 20:24]
  wire  host_dpi_dpi_req_opcode; // @[SimShell.scala 20:24]
  wire [31:0] host_dpi_dpi_req_addr; // @[SimShell.scala 20:24]
  wire [31:0] host_dpi_dpi_req_value; // @[SimShell.scala 20:24]
  wire  host_dpi_dpi_req_deq; // @[SimShell.scala 20:24]
  wire  host_dpi_dpi_resp_valid; // @[SimShell.scala 20:24]
  wire [31:0] host_dpi_dpi_resp_bits; // @[SimShell.scala 20:24]
  wire  host_axi_clock; // @[SimShell.scala 21:24]
  wire  host_axi_reset; // @[SimShell.scala 21:24]
  wire  host_axi_io_dpi_req_valid; // @[SimShell.scala 21:24]
  wire  host_axi_io_dpi_req_opcode; // @[SimShell.scala 21:24]
  wire [31:0] host_axi_io_dpi_req_addr; // @[SimShell.scala 21:24]
  wire [31:0] host_axi_io_dpi_req_value; // @[SimShell.scala 21:24]
  wire  host_axi_io_dpi_req_deq; // @[SimShell.scala 21:24]
  wire  host_axi_io_dpi_resp_valid; // @[SimShell.scala 21:24]
  wire [31:0] host_axi_io_dpi_resp_bits; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_aw_ready; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_aw_valid; // @[SimShell.scala 21:24]
  wire [31:0] host_axi_io_axi_aw_bits_addr; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_w_ready; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_w_valid; // @[SimShell.scala 21:24]
  wire [63:0] host_axi_io_axi_w_bits_data; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_b_ready; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_b_valid; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_ar_ready; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_ar_valid; // @[SimShell.scala 21:24]
  wire [31:0] host_axi_io_axi_ar_bits_addr; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_r_ready; // @[SimShell.scala 21:24]
  wire  host_axi_io_axi_r_valid; // @[SimShell.scala 21:24]
  wire [63:0] host_axi_io_axi_r_bits_data; // @[SimShell.scala 21:24]
  VTAHostDPI host_dpi ( // @[SimShell.scala 20:24]
    .clock(host_dpi_clock),
    .reset(host_dpi_reset),
    .dpi_req_valid(host_dpi_dpi_req_valid),
    .dpi_req_opcode(host_dpi_dpi_req_opcode),
    .dpi_req_addr(host_dpi_dpi_req_addr),
    .dpi_req_value(host_dpi_dpi_req_value),
    .dpi_req_deq(host_dpi_dpi_req_deq),
    .dpi_resp_valid(host_dpi_dpi_resp_valid),
    .dpi_resp_bits(host_dpi_dpi_resp_bits)
  );
  VTAHostDPIToAXI host_axi ( // @[SimShell.scala 21:24]
    .clock(host_axi_clock),
    .reset(host_axi_reset),
    .io_dpi_req_valid(host_axi_io_dpi_req_valid),
    .io_dpi_req_opcode(host_axi_io_dpi_req_opcode),
    .io_dpi_req_addr(host_axi_io_dpi_req_addr),
    .io_dpi_req_value(host_axi_io_dpi_req_value),
    .io_dpi_req_deq(host_axi_io_dpi_req_deq),
    .io_dpi_resp_valid(host_axi_io_dpi_resp_valid),
    .io_dpi_resp_bits(host_axi_io_dpi_resp_bits),
    .io_axi_aw_ready(host_axi_io_axi_aw_ready),
    .io_axi_aw_valid(host_axi_io_axi_aw_valid),
    .io_axi_aw_bits_addr(host_axi_io_axi_aw_bits_addr),
    .io_axi_w_ready(host_axi_io_axi_w_ready),
    .io_axi_w_valid(host_axi_io_axi_w_valid),
    .io_axi_w_bits_data(host_axi_io_axi_w_bits_data),
    .io_axi_b_ready(host_axi_io_axi_b_ready),
    .io_axi_b_valid(host_axi_io_axi_b_valid),
    .io_axi_ar_ready(host_axi_io_axi_ar_ready),
    .io_axi_ar_valid(host_axi_io_axi_ar_valid),
    .io_axi_ar_bits_addr(host_axi_io_axi_ar_bits_addr),
    .io_axi_r_ready(host_axi_io_axi_r_ready),
    .io_axi_r_valid(host_axi_io_axi_r_valid),
    .io_axi_r_bits_data(host_axi_io_axi_r_bits_data)
  );
  assign io_axi_aw_valid = host_axi_io_axi_aw_valid; // @[SimShell.scala 25:10]
  assign io_axi_aw_bits_addr = host_axi_io_axi_aw_bits_addr; // @[SimShell.scala 25:10]
  assign io_axi_w_valid = host_axi_io_axi_w_valid; // @[SimShell.scala 25:10]
  assign io_axi_w_bits_data = host_axi_io_axi_w_bits_data; // @[SimShell.scala 25:10]
  assign io_axi_b_ready = host_axi_io_axi_b_ready; // @[SimShell.scala 25:10]
  assign io_axi_ar_valid = host_axi_io_axi_ar_valid; // @[SimShell.scala 25:10]
  assign io_axi_ar_bits_addr = host_axi_io_axi_ar_bits_addr; // @[SimShell.scala 25:10]
  assign io_axi_r_ready = host_axi_io_axi_r_ready; // @[SimShell.scala 25:10]
  assign host_dpi_clock = clock; // @[SimShell.scala 23:21]
  assign host_dpi_reset = reset; // @[SimShell.scala 22:21]
  assign host_dpi_dpi_req_deq = host_axi_io_dpi_req_deq; // @[SimShell.scala 24:19]
  assign host_dpi_dpi_resp_valid = host_axi_io_dpi_resp_valid; // @[SimShell.scala 24:19]
  assign host_dpi_dpi_resp_bits = host_axi_io_dpi_resp_bits; // @[SimShell.scala 24:19]
  assign host_axi_clock = clock;
  assign host_axi_reset = reset;
  assign host_axi_io_dpi_req_valid = host_dpi_dpi_req_valid; // @[SimShell.scala 24:19]
  assign host_axi_io_dpi_req_opcode = host_dpi_dpi_req_opcode; // @[SimShell.scala 24:19]
  assign host_axi_io_dpi_req_addr = host_dpi_dpi_req_addr; // @[SimShell.scala 24:19]
  assign host_axi_io_dpi_req_value = host_dpi_dpi_req_value; // @[SimShell.scala 24:19]
  assign host_axi_io_axi_aw_ready = io_axi_aw_ready; // @[SimShell.scala 25:10]
  assign host_axi_io_axi_w_ready = io_axi_w_ready; // @[SimShell.scala 25:10]
  assign host_axi_io_axi_b_valid = io_axi_b_valid; // @[SimShell.scala 25:10]
  assign host_axi_io_axi_ar_ready = io_axi_ar_ready; // @[SimShell.scala 25:10]
  assign host_axi_io_axi_r_valid = io_axi_r_valid; // @[SimShell.scala 25:10]
  assign host_axi_io_axi_r_bits_data = io_axi_r_bits_data; // @[SimShell.scala 25:10]
endmodule
module VTAMemDPIToAXI(
  input         clock,
  input         reset,
  output        io_dpi_req_valid,
  output        io_dpi_req_opcode,
  output [31:0] io_dpi_req_len,
  output [63:0] io_dpi_req_addr,
  output        io_dpi_wr_valid,
  output [63:0] io_dpi_wr_bits,
  output        io_dpi_rd_ready,
  input         io_dpi_rd_valid,
  input  [63:0] io_dpi_rd_bits,
  output        io_axi_aw_ready,
  input         io_axi_aw_valid,
  input  [31:0] io_axi_aw_bits_addr,
  input  [31:0] io_axi_aw_bits_len,
  output        io_axi_w_ready,
  input         io_axi_w_valid,
  input  [63:0] io_axi_w_bits_data,
  input         io_axi_w_bits_last,
  input         io_axi_b_ready,
  output        io_axi_b_valid,
  output        io_axi_ar_ready,
  input         io_axi_ar_valid,
  input  [31:0] io_axi_ar_bits_addr,
  input  [31:0] io_axi_ar_bits_len,
  input         io_axi_r_ready,
  output        io_axi_r_valid,
  output [63:0] io_axi_r_bits_data,
  output        io_axi_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  opcode; // @[VTAMemDPI.scala 85:23]
  reg [31:0] len; // @[VTAMemDPI.scala 86:20]
  reg [63:0] addr; // @[VTAMemDPI.scala 87:21]
  reg [2:0] state; // @[VTAMemDPI.scala 90:22]
  wire  _T_2 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = io_axi_r_ready & io_dpi_rd_valid; // @[VTAMemDPI.scala 106:27]
  wire  _T_6 = len == 32'h0; // @[VTAMemDPI.scala 106:53]
  wire  _T_7 = _T_5 & _T_6; // @[VTAMemDPI.scala 106:46]
  wire  _T_8 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_10 = io_axi_w_valid & io_axi_w_bits_last; // @[VTAMemDPI.scala 116:27]
  wire  _T_11 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = state == 3'h0; // @[VTAMemDPI.scala 127:14]
  wire  _GEN_13 = io_axi_aw_valid | opcode; // @[VTAMemDPI.scala 132:33]
  wire  _T_13 = state == 3'h2; // @[VTAMemDPI.scala 138:20]
  wire  _T_15 = len != 32'h0; // @[VTAMemDPI.scala 139:51]
  wire  _T_16 = _T_5 & _T_15; // @[VTAMemDPI.scala 139:44]
  wire [31:0] _T_18 = len - 32'h1; // @[VTAMemDPI.scala 140:18]
  wire  _T_19 = state == 3'h1; // @[VTAMemDPI.scala 144:30]
  wire  _T_20 = _T_19 & io_axi_ar_valid; // @[VTAMemDPI.scala 144:47]
  wire  _T_21 = state == 3'h3; // @[VTAMemDPI.scala 144:75]
  wire  _T_22 = _T_21 & io_axi_aw_valid; // @[VTAMemDPI.scala 144:93]
  wire  _T_31 = state == 3'h4; // @[VTAMemDPI.scala 160:28]
  assign io_dpi_req_valid = _T_20 | _T_22; // @[VTAMemDPI.scala 144:20]
  assign io_dpi_req_opcode = opcode; // @[VTAMemDPI.scala 145:21]
  assign io_dpi_req_len = len; // @[VTAMemDPI.scala 146:18]
  assign io_dpi_req_addr = addr; // @[VTAMemDPI.scala 147:19]
  assign io_dpi_wr_valid = _T_31 & io_axi_w_valid; // @[VTAMemDPI.scala 160:19]
  assign io_dpi_wr_bits = io_axi_w_bits_data; // @[VTAMemDPI.scala 161:18]
  assign io_dpi_rd_ready = _T_13 & io_axi_r_ready; // @[VTAMemDPI.scala 158:19]
  assign io_axi_aw_ready = state == 3'h3; // @[VTAMemDPI.scala 150:19]
  assign io_axi_w_ready = state == 3'h4; // @[VTAMemDPI.scala 162:18]
  assign io_axi_b_valid = state == 3'h5; // @[VTAMemDPI.scala 164:18]
  assign io_axi_ar_ready = state == 3'h1; // @[VTAMemDPI.scala 149:19]
  assign io_axi_r_valid = _T_13 & io_dpi_rd_valid; // @[VTAMemDPI.scala 152:18]
  assign io_axi_r_bits_data = io_dpi_rd_bits; // @[VTAMemDPI.scala 153:22]
  assign io_axi_r_bits_last = len == 32'h0; // @[VTAMemDPI.scala 154:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  opcode = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  len = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  addr = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      opcode <= 1'h0;
    end else if (_T_12) begin
      if (io_axi_ar_valid) begin
        opcode <= 1'h0;
      end else begin
        opcode <= _GEN_13;
      end
    end
    if (reset) begin
      len <= 32'h0;
    end else if (_T_12) begin
      if (io_axi_ar_valid) begin
        len <= io_axi_ar_bits_len;
      end else if (io_axi_aw_valid) begin
        len <= io_axi_aw_bits_len;
      end
    end else if (_T_13) begin
      if (_T_16) begin
        len <= _T_18;
      end
    end
    if (reset) begin
      addr <= 64'h0;
    end else if (_T_12) begin
      if (io_axi_ar_valid) begin
        addr <= {{32'd0}, io_axi_ar_bits_addr};
      end else if (io_axi_aw_valid) begin
        addr <= {{32'd0}, io_axi_aw_bits_addr};
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_2) begin
      if (io_axi_ar_valid) begin
        state <= 3'h1;
      end else if (io_axi_aw_valid) begin
        state <= 3'h3;
      end
    end else if (_T_3) begin
      if (io_axi_ar_valid) begin
        state <= 3'h2;
      end
    end else if (_T_4) begin
      if (_T_7) begin
        state <= 3'h0;
      end
    end else if (_T_8) begin
      if (io_axi_aw_valid) begin
        state <= 3'h4;
      end
    end else if (_T_9) begin
      if (_T_10) begin
        state <= 3'h5;
      end
    end else if (_T_11) begin
      if (io_axi_b_ready) begin
        state <= 3'h0;
      end
    end
  end
endmodule
module VTAMem(
  input         clock,
  input         reset,
  output        io_axi_aw_ready,
  input         io_axi_aw_valid,
  input  [31:0] io_axi_aw_bits_addr,
  input  [31:0] io_axi_aw_bits_len,
  output        io_axi_w_ready,
  input         io_axi_w_valid,
  input  [63:0] io_axi_w_bits_data,
  input         io_axi_w_bits_last,
  input         io_axi_b_ready,
  output        io_axi_b_valid,
  output        io_axi_ar_ready,
  input         io_axi_ar_valid,
  input  [31:0] io_axi_ar_bits_addr,
  input  [31:0] io_axi_ar_bits_len,
  input         io_axi_r_ready,
  output        io_axi_r_valid,
  output [63:0] io_axi_r_bits_data,
  output        io_axi_r_bits_last
);
  wire  mem_dpi_clock; // @[SimShell.scala 38:23]
  wire  mem_dpi_reset; // @[SimShell.scala 38:23]
  wire  mem_dpi_dpi_req_valid; // @[SimShell.scala 38:23]
  wire  mem_dpi_dpi_req_opcode; // @[SimShell.scala 38:23]
  wire [31:0] mem_dpi_dpi_req_len; // @[SimShell.scala 38:23]
  wire [63:0] mem_dpi_dpi_req_addr; // @[SimShell.scala 38:23]
  wire  mem_dpi_dpi_wr_valid; // @[SimShell.scala 38:23]
  wire [63:0] mem_dpi_dpi_wr_bits; // @[SimShell.scala 38:23]
  wire  mem_dpi_dpi_rd_ready; // @[SimShell.scala 38:23]
  wire  mem_dpi_dpi_rd_valid; // @[SimShell.scala 38:23]
  wire [63:0] mem_dpi_dpi_rd_bits; // @[SimShell.scala 38:23]
  wire  mem_axi_clock; // @[SimShell.scala 39:23]
  wire  mem_axi_reset; // @[SimShell.scala 39:23]
  wire  mem_axi_io_dpi_req_valid; // @[SimShell.scala 39:23]
  wire  mem_axi_io_dpi_req_opcode; // @[SimShell.scala 39:23]
  wire [31:0] mem_axi_io_dpi_req_len; // @[SimShell.scala 39:23]
  wire [63:0] mem_axi_io_dpi_req_addr; // @[SimShell.scala 39:23]
  wire  mem_axi_io_dpi_wr_valid; // @[SimShell.scala 39:23]
  wire [63:0] mem_axi_io_dpi_wr_bits; // @[SimShell.scala 39:23]
  wire  mem_axi_io_dpi_rd_ready; // @[SimShell.scala 39:23]
  wire  mem_axi_io_dpi_rd_valid; // @[SimShell.scala 39:23]
  wire [63:0] mem_axi_io_dpi_rd_bits; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_aw_ready; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_aw_valid; // @[SimShell.scala 39:23]
  wire [31:0] mem_axi_io_axi_aw_bits_addr; // @[SimShell.scala 39:23]
  wire [31:0] mem_axi_io_axi_aw_bits_len; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_w_ready; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_w_valid; // @[SimShell.scala 39:23]
  wire [63:0] mem_axi_io_axi_w_bits_data; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_w_bits_last; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_b_ready; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_b_valid; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_ar_ready; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_ar_valid; // @[SimShell.scala 39:23]
  wire [31:0] mem_axi_io_axi_ar_bits_addr; // @[SimShell.scala 39:23]
  wire [31:0] mem_axi_io_axi_ar_bits_len; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_r_ready; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_r_valid; // @[SimShell.scala 39:23]
  wire [63:0] mem_axi_io_axi_r_bits_data; // @[SimShell.scala 39:23]
  wire  mem_axi_io_axi_r_bits_last; // @[SimShell.scala 39:23]
  VTAMemDPI mem_dpi ( // @[SimShell.scala 38:23]
    .clock(mem_dpi_clock),
    .reset(mem_dpi_reset),
    .dpi_req_valid(mem_dpi_dpi_req_valid),
    .dpi_req_opcode(mem_dpi_dpi_req_opcode),
    .dpi_req_len(mem_dpi_dpi_req_len),
    .dpi_req_addr(mem_dpi_dpi_req_addr),
    .dpi_wr_valid(mem_dpi_dpi_wr_valid),
    .dpi_wr_bits(mem_dpi_dpi_wr_bits),
    .dpi_rd_ready(mem_dpi_dpi_rd_ready),
    .dpi_rd_valid(mem_dpi_dpi_rd_valid),
    .dpi_rd_bits(mem_dpi_dpi_rd_bits)
  );
  VTAMemDPIToAXI mem_axi ( // @[SimShell.scala 39:23]
    .clock(mem_axi_clock),
    .reset(mem_axi_reset),
    .io_dpi_req_valid(mem_axi_io_dpi_req_valid),
    .io_dpi_req_opcode(mem_axi_io_dpi_req_opcode),
    .io_dpi_req_len(mem_axi_io_dpi_req_len),
    .io_dpi_req_addr(mem_axi_io_dpi_req_addr),
    .io_dpi_wr_valid(mem_axi_io_dpi_wr_valid),
    .io_dpi_wr_bits(mem_axi_io_dpi_wr_bits),
    .io_dpi_rd_ready(mem_axi_io_dpi_rd_ready),
    .io_dpi_rd_valid(mem_axi_io_dpi_rd_valid),
    .io_dpi_rd_bits(mem_axi_io_dpi_rd_bits),
    .io_axi_aw_ready(mem_axi_io_axi_aw_ready),
    .io_axi_aw_valid(mem_axi_io_axi_aw_valid),
    .io_axi_aw_bits_addr(mem_axi_io_axi_aw_bits_addr),
    .io_axi_aw_bits_len(mem_axi_io_axi_aw_bits_len),
    .io_axi_w_ready(mem_axi_io_axi_w_ready),
    .io_axi_w_valid(mem_axi_io_axi_w_valid),
    .io_axi_w_bits_data(mem_axi_io_axi_w_bits_data),
    .io_axi_w_bits_last(mem_axi_io_axi_w_bits_last),
    .io_axi_b_ready(mem_axi_io_axi_b_ready),
    .io_axi_b_valid(mem_axi_io_axi_b_valid),
    .io_axi_ar_ready(mem_axi_io_axi_ar_ready),
    .io_axi_ar_valid(mem_axi_io_axi_ar_valid),
    .io_axi_ar_bits_addr(mem_axi_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(mem_axi_io_axi_ar_bits_len),
    .io_axi_r_ready(mem_axi_io_axi_r_ready),
    .io_axi_r_valid(mem_axi_io_axi_r_valid),
    .io_axi_r_bits_data(mem_axi_io_axi_r_bits_data),
    .io_axi_r_bits_last(mem_axi_io_axi_r_bits_last)
  );
  assign io_axi_aw_ready = mem_axi_io_axi_aw_ready; // @[SimShell.scala 43:10]
  assign io_axi_w_ready = mem_axi_io_axi_w_ready; // @[SimShell.scala 43:10]
  assign io_axi_b_valid = mem_axi_io_axi_b_valid; // @[SimShell.scala 43:10]
  assign io_axi_ar_ready = mem_axi_io_axi_ar_ready; // @[SimShell.scala 43:10]
  assign io_axi_r_valid = mem_axi_io_axi_r_valid; // @[SimShell.scala 43:10]
  assign io_axi_r_bits_data = mem_axi_io_axi_r_bits_data; // @[SimShell.scala 43:10]
  assign io_axi_r_bits_last = mem_axi_io_axi_r_bits_last; // @[SimShell.scala 43:10]
  assign mem_dpi_clock = clock; // @[SimShell.scala 41:20]
  assign mem_dpi_reset = reset; // @[SimShell.scala 40:20]
  assign mem_dpi_dpi_req_valid = mem_axi_io_dpi_req_valid; // @[SimShell.scala 42:18]
  assign mem_dpi_dpi_req_opcode = mem_axi_io_dpi_req_opcode; // @[SimShell.scala 42:18]
  assign mem_dpi_dpi_req_len = mem_axi_io_dpi_req_len; // @[SimShell.scala 42:18]
  assign mem_dpi_dpi_req_addr = mem_axi_io_dpi_req_addr; // @[SimShell.scala 42:18]
  assign mem_dpi_dpi_wr_valid = mem_axi_io_dpi_wr_valid; // @[SimShell.scala 42:18]
  assign mem_dpi_dpi_wr_bits = mem_axi_io_dpi_wr_bits; // @[SimShell.scala 42:18]
  assign mem_dpi_dpi_rd_ready = mem_axi_io_dpi_rd_ready; // @[SimShell.scala 42:18]
  assign mem_axi_clock = clock;
  assign mem_axi_reset = reset;
  assign mem_axi_io_dpi_rd_valid = mem_dpi_dpi_rd_valid; // @[SimShell.scala 42:18]
  assign mem_axi_io_dpi_rd_bits = mem_dpi_dpi_rd_bits; // @[SimShell.scala 42:18]
  assign mem_axi_io_axi_aw_valid = io_axi_aw_valid; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_aw_bits_addr = io_axi_aw_bits_addr; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_aw_bits_len = io_axi_aw_bits_len; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_w_valid = io_axi_w_valid; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_w_bits_data = io_axi_w_bits_data; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_w_bits_last = io_axi_w_bits_last; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_b_ready = io_axi_b_ready; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_ar_valid = io_axi_ar_valid; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_ar_bits_addr = io_axi_ar_bits_addr; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_ar_bits_len = io_axi_ar_bits_len; // @[SimShell.scala 43:10]
  assign mem_axi_io_axi_r_ready = io_axi_r_ready; // @[SimShell.scala 43:10]
endmodule
module AXISimShell(
  input         clock,
  input         reset,
  output        mem_aw_ready,
  input         mem_aw_valid,
  input  [31:0] mem_aw_bits_addr,
  input  [31:0] mem_aw_bits_len,
  output        mem_w_ready,
  input         mem_w_valid,
  input  [63:0] mem_w_bits_data,
  input         mem_w_bits_last,
  input         mem_b_ready,
  output        mem_b_valid,
  output        mem_ar_ready,
  input         mem_ar_valid,
  input  [31:0] mem_ar_bits_addr,
  input  [31:0] mem_ar_bits_len,
  input         mem_r_ready,
  output        mem_r_valid,
  output [63:0] mem_r_bits_data,
  output        mem_r_bits_last,
  input         host_aw_ready,
  output        host_aw_valid,
  output [31:0] host_aw_bits_addr,
  input         host_w_ready,
  output        host_w_valid,
  output [63:0] host_w_bits_data,
  output        host_b_ready,
  input         host_b_valid,
  input         host_ar_ready,
  output        host_ar_valid,
  output [31:0] host_ar_bits_addr,
  output        host_r_ready,
  input         host_r_valid,
  input  [63:0] host_r_bits_data,
  input         sim_clock,
  output        sim_wait
);
  wire  mod_sim_clock; // @[SimShell.scala 93:23]
  wire  mod_sim_reset; // @[SimShell.scala 93:23]
  wire  mod_sim_sim_wait; // @[SimShell.scala 93:23]
  wire  mod_host_clock; // @[SimShell.scala 94:24]
  wire  mod_host_reset; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_aw_ready; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_aw_valid; // @[SimShell.scala 94:24]
  wire [31:0] mod_host_io_axi_aw_bits_addr; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_w_ready; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_w_valid; // @[SimShell.scala 94:24]
  wire [63:0] mod_host_io_axi_w_bits_data; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_b_ready; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_b_valid; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_ar_ready; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_ar_valid; // @[SimShell.scala 94:24]
  wire [31:0] mod_host_io_axi_ar_bits_addr; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_r_ready; // @[SimShell.scala 94:24]
  wire  mod_host_io_axi_r_valid; // @[SimShell.scala 94:24]
  wire [63:0] mod_host_io_axi_r_bits_data; // @[SimShell.scala 94:24]
  wire  mod_mem_clock; // @[SimShell.scala 95:23]
  wire  mod_mem_reset; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_aw_ready; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_aw_valid; // @[SimShell.scala 95:23]
  wire [31:0] mod_mem_io_axi_aw_bits_addr; // @[SimShell.scala 95:23]
  wire [31:0] mod_mem_io_axi_aw_bits_len; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_w_ready; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_w_valid; // @[SimShell.scala 95:23]
  wire [63:0] mod_mem_io_axi_w_bits_data; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_w_bits_last; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_b_ready; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_b_valid; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_ar_ready; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_ar_valid; // @[SimShell.scala 95:23]
  wire [31:0] mod_mem_io_axi_ar_bits_addr; // @[SimShell.scala 95:23]
  wire [31:0] mod_mem_io_axi_ar_bits_len; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_r_ready; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_r_valid; // @[SimShell.scala 95:23]
  wire [63:0] mod_mem_io_axi_r_bits_data; // @[SimShell.scala 95:23]
  wire  mod_mem_io_axi_r_bits_last; // @[SimShell.scala 95:23]
  VTASim mod_sim ( // @[SimShell.scala 93:23]
    .clock(mod_sim_clock),
    .reset(mod_sim_reset),
    .sim_wait(mod_sim_sim_wait)
  );
  VTAHost mod_host ( // @[SimShell.scala 94:24]
    .clock(mod_host_clock),
    .reset(mod_host_reset),
    .io_axi_aw_ready(mod_host_io_axi_aw_ready),
    .io_axi_aw_valid(mod_host_io_axi_aw_valid),
    .io_axi_aw_bits_addr(mod_host_io_axi_aw_bits_addr),
    .io_axi_w_ready(mod_host_io_axi_w_ready),
    .io_axi_w_valid(mod_host_io_axi_w_valid),
    .io_axi_w_bits_data(mod_host_io_axi_w_bits_data),
    .io_axi_b_ready(mod_host_io_axi_b_ready),
    .io_axi_b_valid(mod_host_io_axi_b_valid),
    .io_axi_ar_ready(mod_host_io_axi_ar_ready),
    .io_axi_ar_valid(mod_host_io_axi_ar_valid),
    .io_axi_ar_bits_addr(mod_host_io_axi_ar_bits_addr),
    .io_axi_r_ready(mod_host_io_axi_r_ready),
    .io_axi_r_valid(mod_host_io_axi_r_valid),
    .io_axi_r_bits_data(mod_host_io_axi_r_bits_data)
  );
  VTAMem mod_mem ( // @[SimShell.scala 95:23]
    .clock(mod_mem_clock),
    .reset(mod_mem_reset),
    .io_axi_aw_ready(mod_mem_io_axi_aw_ready),
    .io_axi_aw_valid(mod_mem_io_axi_aw_valid),
    .io_axi_aw_bits_addr(mod_mem_io_axi_aw_bits_addr),
    .io_axi_aw_bits_len(mod_mem_io_axi_aw_bits_len),
    .io_axi_w_ready(mod_mem_io_axi_w_ready),
    .io_axi_w_valid(mod_mem_io_axi_w_valid),
    .io_axi_w_bits_data(mod_mem_io_axi_w_bits_data),
    .io_axi_w_bits_last(mod_mem_io_axi_w_bits_last),
    .io_axi_b_ready(mod_mem_io_axi_b_ready),
    .io_axi_b_valid(mod_mem_io_axi_b_valid),
    .io_axi_ar_ready(mod_mem_io_axi_ar_ready),
    .io_axi_ar_valid(mod_mem_io_axi_ar_valid),
    .io_axi_ar_bits_addr(mod_mem_io_axi_ar_bits_addr),
    .io_axi_ar_bits_len(mod_mem_io_axi_ar_bits_len),
    .io_axi_r_ready(mod_mem_io_axi_r_ready),
    .io_axi_r_valid(mod_mem_io_axi_r_valid),
    .io_axi_r_bits_data(mod_mem_io_axi_r_bits_data),
    .io_axi_r_bits_last(mod_mem_io_axi_r_bits_last)
  );
  assign mem_aw_ready = mod_mem_io_axi_aw_ready; // @[SimShell.scala 96:7]
  assign mem_w_ready = mod_mem_io_axi_w_ready; // @[SimShell.scala 96:7]
  assign mem_b_valid = mod_mem_io_axi_b_valid; // @[SimShell.scala 96:7]
  assign mem_ar_ready = mod_mem_io_axi_ar_ready; // @[SimShell.scala 96:7]
  assign mem_r_valid = mod_mem_io_axi_r_valid; // @[SimShell.scala 96:7]
  assign mem_r_bits_data = mod_mem_io_axi_r_bits_data; // @[SimShell.scala 96:7]
  assign mem_r_bits_last = mod_mem_io_axi_r_bits_last; // @[SimShell.scala 96:7]
  assign host_aw_valid = mod_host_io_axi_aw_valid; // @[SimShell.scala 97:8]
  assign host_aw_bits_addr = mod_host_io_axi_aw_bits_addr; // @[SimShell.scala 97:8]
  assign host_w_valid = mod_host_io_axi_w_valid; // @[SimShell.scala 97:8]
  assign host_w_bits_data = mod_host_io_axi_w_bits_data; // @[SimShell.scala 97:8]
  assign host_b_ready = mod_host_io_axi_b_ready; // @[SimShell.scala 97:8]
  assign host_ar_valid = mod_host_io_axi_ar_valid; // @[SimShell.scala 97:8]
  assign host_ar_bits_addr = mod_host_io_axi_ar_bits_addr; // @[SimShell.scala 97:8]
  assign host_r_ready = mod_host_io_axi_r_ready; // @[SimShell.scala 97:8]
  assign sim_wait = mod_sim_sim_wait; // @[SimShell.scala 100:12]
  assign mod_sim_clock = sim_clock; // @[SimShell.scala 99:17]
  assign mod_sim_reset = reset; // @[SimShell.scala 98:17]
  assign mod_host_clock = clock;
  assign mod_host_reset = reset;
  assign mod_host_io_axi_aw_ready = host_aw_ready; // @[SimShell.scala 97:8]
  assign mod_host_io_axi_w_ready = host_w_ready; // @[SimShell.scala 97:8]
  assign mod_host_io_axi_b_valid = host_b_valid; // @[SimShell.scala 97:8]
  assign mod_host_io_axi_ar_ready = host_ar_ready; // @[SimShell.scala 97:8]
  assign mod_host_io_axi_r_valid = host_r_valid; // @[SimShell.scala 97:8]
  assign mod_host_io_axi_r_bits_data = host_r_bits_data; // @[SimShell.scala 97:8]
  assign mod_mem_clock = clock;
  assign mod_mem_reset = reset;
  assign mod_mem_io_axi_aw_valid = mem_aw_valid; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_aw_bits_addr = mem_aw_bits_addr; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_aw_bits_len = mem_aw_bits_len; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_w_valid = mem_w_valid; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_w_bits_data = mem_w_bits_data; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_w_bits_last = mem_w_bits_last; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_b_ready = mem_b_ready; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_ar_valid = mem_ar_valid; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_ar_bits_addr = mem_ar_bits_addr; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_ar_bits_len = mem_ar_bits_len; // @[SimShell.scala 96:7]
  assign mod_mem_io_axi_r_ready = mem_r_ready; // @[SimShell.scala 96:7]
endmodule
module DCR(
  input         clock,
  input         reset,
  output        io_host_aw_ready,
  input         io_host_aw_valid,
  input  [31:0] io_host_aw_bits_addr,
  output        io_host_w_ready,
  input         io_host_w_valid,
  input  [63:0] io_host_w_bits_data,
  input         io_host_b_ready,
  output        io_host_b_valid,
  output        io_host_ar_ready,
  input         io_host_ar_valid,
  input  [31:0] io_host_ar_bits_addr,
  input         io_host_r_ready,
  output        io_host_r_valid,
  output [63:0] io_host_r_bits_data,
  output        io_dcr_launch,
  input         io_dcr_finish,
  input         io_dcr_ecnt_0_valid,
  input  [31:0] io_dcr_ecnt_0_bits,
  input  [31:0] io_dcr_ecnt_1_bits,
  input  [31:0] io_dcr_ecnt_2_bits,
  input  [31:0] io_dcr_ecnt_3_bits,
  input  [31:0] io_dcr_ecnt_4_bits,
  input  [31:0] io_dcr_ecnt_5_bits,
  input  [31:0] io_dcr_ecnt_6_bits,
  output [31:0] io_dcr_vals_0,
  output [31:0] io_dcr_ptrs_1,
  output [31:0] io_dcr_ptrs_2,
  output [31:0] io_dcr_ptrs_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] waddr; // @[DCR.scala 88:22]
  reg [1:0] wstate; // @[DCR.scala 91:23]
  reg  rstate; // @[DCR.scala 95:23]
  reg [31:0] rdata; // @[DCR.scala 96:22]
  reg [31:0] reg_0; // @[DCR.scala 102:37]
  reg [31:0] reg_1; // @[DCR.scala 102:37]
  reg [31:0] reg_2; // @[DCR.scala 102:37]
  reg [31:0] reg_3; // @[DCR.scala 102:37]
  reg [31:0] reg_4; // @[DCR.scala 102:37]
  reg [31:0] reg_5; // @[DCR.scala 102:37]
  reg [31:0] reg_6; // @[DCR.scala 102:37]
  reg [31:0] reg_7; // @[DCR.scala 102:37]
  reg [31:0] reg_18; // @[DCR.scala 102:37]
  reg [31:0] reg_19; // @[DCR.scala 102:37]
  reg [31:0] reg_20; // @[DCR.scala 102:37]
  reg [31:0] reg_21; // @[DCR.scala 102:37]
  reg [31:0] reg_22; // @[DCR.scala 102:37]
  wire  _T = 2'h0 == wstate; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == wstate; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h2 == wstate; // @[Conditional.scala 37:30]
  wire  _T_3 = io_host_aw_ready & io_host_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_7 = ~rstate; // @[Conditional.scala 37:30]
  wire  _GEN_7 = io_host_ar_valid | rstate; // @[DCR.scala 138:30]
  wire  _T_11 = io_host_w_ready & io_host_w_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = 32'h0 == waddr; // @[DCR.scala 156:44]
  wire  _T_13 = _T_11 & _T_12; // @[DCR.scala 156:31]
  wire [63:0] _GEN_11 = _T_13 ? io_host_w_bits_data : {{32'd0}, reg_0}; // @[DCR.scala 156:55]
  wire [63:0] _GEN_12 = io_dcr_finish ? 64'h2 : _GEN_11; // @[DCR.scala 154:23]
  wire  _T_15 = 32'h4 == waddr; // @[DCR.scala 163:51]
  wire  _T_16 = _T_11 & _T_15; // @[DCR.scala 163:33]
  wire [63:0] _GEN_13 = _T_16 ? io_host_w_bits_data : {{32'd0}, reg_1}; // @[DCR.scala 163:62]
  wire [63:0] _GEN_14 = io_dcr_ecnt_0_valid ? {{32'd0}, io_dcr_ecnt_0_bits} : _GEN_13; // @[DCR.scala 161:32]
  wire [63:0] _GEN_16 = {{32'd0}, io_dcr_ecnt_1_bits}; // @[DCR.scala 161:32]
  wire [63:0] _GEN_18 = {{32'd0}, io_dcr_ecnt_2_bits}; // @[DCR.scala 161:32]
  wire [63:0] _GEN_20 = {{32'd0}, io_dcr_ecnt_3_bits}; // @[DCR.scala 161:32]
  wire [63:0] _GEN_22 = {{32'd0}, io_dcr_ecnt_4_bits}; // @[DCR.scala 161:32]
  wire [63:0] _GEN_24 = {{32'd0}, io_dcr_ecnt_5_bits}; // @[DCR.scala 161:32]
  wire [63:0] _GEN_26 = {{32'd0}, io_dcr_ecnt_6_bits}; // @[DCR.scala 161:32]
  wire  _T_66 = 32'h48 == waddr; // @[DCR.scala 169:45]
  wire  _T_67 = _T_11 & _T_66; // @[DCR.scala 169:27]
  wire [63:0] _GEN_47 = _T_67 ? io_host_w_bits_data : {{32'd0}, reg_18}; // @[DCR.scala 169:56]
  wire  _T_69 = 32'h4c == waddr; // @[DCR.scala 169:45]
  wire  _T_70 = _T_11 & _T_69; // @[DCR.scala 169:27]
  wire [63:0] _GEN_48 = _T_70 ? io_host_w_bits_data : {{32'd0}, reg_19}; // @[DCR.scala 169:56]
  wire  _T_72 = 32'h50 == waddr; // @[DCR.scala 169:45]
  wire  _T_73 = _T_11 & _T_72; // @[DCR.scala 169:27]
  wire [63:0] _GEN_49 = _T_73 ? io_host_w_bits_data : {{32'd0}, reg_20}; // @[DCR.scala 169:56]
  wire  _T_75 = 32'h54 == waddr; // @[DCR.scala 169:45]
  wire  _T_76 = _T_11 & _T_75; // @[DCR.scala 169:27]
  wire [63:0] _GEN_50 = _T_76 ? io_host_w_bits_data : {{32'd0}, reg_21}; // @[DCR.scala 169:56]
  wire  _T_78 = 32'h58 == waddr; // @[DCR.scala 169:45]
  wire  _T_79 = _T_11 & _T_78; // @[DCR.scala 169:27]
  wire [63:0] _GEN_51 = _T_79 ? io_host_w_bits_data : {{32'd0}, reg_22}; // @[DCR.scala 169:56]
  wire  _T_80 = io_host_ar_ready & io_host_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_81 = 32'h0 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_83 = 32'h4 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_85 = 32'h8 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_87 = 32'hc == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_89 = 32'h10 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_91 = 32'h14 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_93 = 32'h18 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_95 = 32'h1c == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_97 = 32'h20 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_99 = 32'h24 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_101 = 32'h28 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_103 = 32'h2c == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_105 = 32'h30 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_107 = 32'h34 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_109 = 32'h38 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_111 = 32'h3c == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_113 = 32'h40 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_115 = 32'h44 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_117 = 32'h48 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_119 = 32'h4c == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_121 = 32'h50 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_123 = 32'h54 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_125 = 32'h58 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  assign io_host_aw_ready = wstate == 2'h0; // @[DCR.scala 131:20]
  assign io_host_w_ready = wstate == 2'h1; // @[DCR.scala 132:19]
  assign io_host_b_valid = wstate == 2'h2; // @[DCR.scala 133:19]
  assign io_host_ar_ready = ~rstate; // @[DCR.scala 149:20]
  assign io_host_r_valid = rstate; // @[DCR.scala 150:19]
  assign io_host_r_bits_data = {{32'd0}, rdata}; // @[DCR.scala 151:23]
  assign io_dcr_launch = reg_0[0]; // @[DCR.scala 178:17]
  assign io_dcr_vals_0 = reg_18; // @[DCR.scala 181:20]
  assign io_dcr_ptrs_1 = reg_20; // @[DCR.scala 186:22]
  assign io_dcr_ptrs_2 = reg_21; // @[DCR.scala 186:22]
  assign io_dcr_ptrs_3 = reg_22; // @[DCR.scala 186:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waddr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  wstate = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  rstate = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  rdata = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_0 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_4 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_5 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_6 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_7 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_18 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_19 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_20 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_21 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_22 = _RAND_16[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      waddr <= 32'hffff;
    end else if (_T_3) begin
      waddr <= io_host_aw_bits_addr;
    end
    if (reset) begin
      wstate <= 2'h0;
    end else if (_T) begin
      if (io_host_aw_valid) begin
        wstate <= 2'h1;
      end
    end else if (_T_1) begin
      if (io_host_w_valid) begin
        wstate <= 2'h2;
      end
    end else if (_T_2) begin
      if (io_host_b_ready) begin
        wstate <= 2'h0;
      end
    end
    if (reset) begin
      rstate <= 1'h0;
    end else if (_T_7) begin
      rstate <= _GEN_7;
    end else if (rstate) begin
      if (io_host_r_ready) begin
        rstate <= 1'h0;
      end
    end
    if (reset) begin
      rdata <= 32'h0;
    end else if (_T_80) begin
      if (_T_125) begin
        rdata <= reg_22;
      end else if (_T_123) begin
        rdata <= reg_21;
      end else if (_T_121) begin
        rdata <= reg_20;
      end else if (_T_119) begin
        rdata <= reg_19;
      end else if (_T_117) begin
        rdata <= reg_18;
      end else if (_T_115) begin
        rdata <= 32'h0;
      end else if (_T_113) begin
        rdata <= 32'h0;
      end else if (_T_111) begin
        rdata <= 32'h0;
      end else if (_T_109) begin
        rdata <= 32'h0;
      end else if (_T_107) begin
        rdata <= 32'h0;
      end else if (_T_105) begin
        rdata <= 32'h0;
      end else if (_T_103) begin
        rdata <= 32'h0;
      end else if (_T_101) begin
        rdata <= 32'h0;
      end else if (_T_99) begin
        rdata <= 32'h0;
      end else if (_T_97) begin
        rdata <= 32'h0;
      end else if (_T_95) begin
        rdata <= reg_7;
      end else if (_T_93) begin
        rdata <= reg_6;
      end else if (_T_91) begin
        rdata <= reg_5;
      end else if (_T_89) begin
        rdata <= reg_4;
      end else if (_T_87) begin
        rdata <= reg_3;
      end else if (_T_85) begin
        rdata <= reg_2;
      end else if (_T_83) begin
        rdata <= reg_1;
      end else if (_T_81) begin
        rdata <= reg_0;
      end else begin
        rdata <= 32'h0;
      end
    end
    if (reset) begin
      reg_0 <= 32'h0;
    end else begin
      reg_0 <= _GEN_12[31:0];
    end
    if (reset) begin
      reg_1 <= 32'h0;
    end else begin
      reg_1 <= _GEN_14[31:0];
    end
    if (reset) begin
      reg_2 <= 32'h0;
    end else begin
      reg_2 <= _GEN_16[31:0];
    end
    if (reset) begin
      reg_3 <= 32'h0;
    end else begin
      reg_3 <= _GEN_18[31:0];
    end
    if (reset) begin
      reg_4 <= 32'h0;
    end else begin
      reg_4 <= _GEN_20[31:0];
    end
    if (reset) begin
      reg_5 <= 32'h0;
    end else begin
      reg_5 <= _GEN_22[31:0];
    end
    if (reset) begin
      reg_6 <= 32'h0;
    end else begin
      reg_6 <= _GEN_24[31:0];
    end
    if (reset) begin
      reg_7 <= 32'h0;
    end else begin
      reg_7 <= _GEN_26[31:0];
    end
    if (reset) begin
      reg_18 <= 32'h0;
    end else begin
      reg_18 <= _GEN_47[31:0];
    end
    if (reset) begin
      reg_19 <= 32'h0;
    end else begin
      reg_19 <= _GEN_48[31:0];
    end
    if (reset) begin
      reg_20 <= 32'h0;
    end else begin
      reg_20 <= _GEN_49[31:0];
    end
    if (reset) begin
      reg_21 <= 32'h0;
    end else begin
      reg_21 <= _GEN_50[31:0];
    end
    if (reset) begin
      reg_22 <= 32'h0;
    end else begin
      reg_22 <= _GEN_51[31:0];
    end
  end
endmodule
module Arbiter(
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [1:0]  io_chosen
);
  wire [1:0] _GEN_0 = io_in_1_valid ? 2'h1 : 2'h2; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_2 = io_in_1_valid ? io_in_1_bits_addr : io_in_2_bits_addr; // @[Arbiter.scala 126:27]
  wire  _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  grant_2 = ~_T; // @[Arbiter.scala 31:78]
  wire  _T_4 = ~grant_2; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_4 | io_in_2_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_2; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_chosen = io_in_0_valid ? 2'h0 : _GEN_0; // @[Arbiter.scala 123:13 Arbiter.scala 127:17 Arbiter.scala 127:17]
endmodule
module DME(
  input         clock,
  input         reset,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output        io_mem_w_bits_last,
  output        io_mem_b_ready,
  input         io_mem_b_valid,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last,
  input         io_dme_rd_0_cmd_valid,
  input  [31:0] io_dme_rd_0_cmd_bits_addr,
  input         io_dme_rd_0_data_ready,
  output        io_dme_rd_0_data_valid,
  output [63:0] io_dme_rd_0_data_bits,
  input         io_dme_rd_1_cmd_valid,
  input  [31:0] io_dme_rd_1_cmd_bits_addr,
  input         io_dme_rd_1_data_ready,
  output        io_dme_rd_1_data_valid,
  output [63:0] io_dme_rd_1_data_bits,
  input         io_dme_rd_2_cmd_valid,
  input  [31:0] io_dme_rd_2_cmd_bits_addr,
  input         io_dme_rd_2_data_ready,
  output        io_dme_rd_2_data_valid,
  output [63:0] io_dme_rd_2_data_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  rd_arb_io_in_0_valid; // @[DME.scala 130:22]
  wire [31:0] rd_arb_io_in_0_bits_addr; // @[DME.scala 130:22]
  wire  rd_arb_io_in_1_valid; // @[DME.scala 130:22]
  wire [31:0] rd_arb_io_in_1_bits_addr; // @[DME.scala 130:22]
  wire  rd_arb_io_in_2_valid; // @[DME.scala 130:22]
  wire [31:0] rd_arb_io_in_2_bits_addr; // @[DME.scala 130:22]
  wire  rd_arb_io_out_ready; // @[DME.scala 130:22]
  wire  rd_arb_io_out_valid; // @[DME.scala 130:22]
  wire [31:0] rd_arb_io_out_bits_addr; // @[DME.scala 130:22]
  wire [1:0] rd_arb_io_chosen; // @[DME.scala 130:22]
  wire  _T = rd_arb_io_out_ready & rd_arb_io_out_valid; // @[Decoupled.scala 40:37]
  reg [1:0] rd_arb_chosen; // @[Reg.scala 15:16]
  reg [1:0] rstate; // @[DME.scala 138:23]
  wire  _T_1 = 2'h0 == rstate; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h1 == rstate; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h2 == rstate; // @[Conditional.scala 37:30]
  wire  _T_4 = io_mem_r_ready & io_mem_r_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = _T_4 & io_mem_r_bits_last; // @[DME.scala 152:28]
  reg [1:0] wstate; // @[DME.scala 168:23]
  reg [31:0] wr_cnt; // @[DME.scala 171:23]
  wire  _T_7 = wstate == 2'h0; // @[DME.scala 174:15]
  wire  _T_8 = io_mem_w_ready & io_mem_w_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _T_10 = wr_cnt + 32'h1; // @[DME.scala 177:22]
  wire  _T_11 = 2'h0 == wstate; // @[Conditional.scala 37:30]
  wire  _T_12 = 2'h1 == wstate; // @[Conditional.scala 37:30]
  wire  _T_13 = 2'h2 == wstate; // @[Conditional.scala 37:30]
  wire  _T_17 = 2'h3 == wstate; // @[Conditional.scala 37:30]
  reg [31:0] rd_addr; // @[Reg.scala 27:20]
  wire  _T_24 = rd_arb_chosen == 2'h0; // @[DME.scala 215:46]
  wire  _T_26 = rd_arb_chosen == 2'h1; // @[DME.scala 215:46]
  wire  _T_28 = rd_arb_chosen == 2'h2; // @[DME.scala 215:46]
  wire  _T_43 = rstate == 2'h2; // @[DME.scala 240:28]
  wire  _GEN_33 = 2'h1 == rd_arb_chosen ? io_dme_rd_1_data_ready : io_dme_rd_0_data_ready; // @[DME.scala 240:42]
  wire  _GEN_40 = 2'h2 == rd_arb_chosen ? io_dme_rd_2_data_ready : _GEN_33; // @[DME.scala 240:42]
  Arbiter rd_arb ( // @[DME.scala 130:22]
    .io_in_0_valid(rd_arb_io_in_0_valid),
    .io_in_0_bits_addr(rd_arb_io_in_0_bits_addr),
    .io_in_1_valid(rd_arb_io_in_1_valid),
    .io_in_1_bits_addr(rd_arb_io_in_1_bits_addr),
    .io_in_2_valid(rd_arb_io_in_2_valid),
    .io_in_2_bits_addr(rd_arb_io_in_2_bits_addr),
    .io_out_ready(rd_arb_io_out_ready),
    .io_out_valid(rd_arb_io_out_valid),
    .io_out_bits_addr(rd_arb_io_out_bits_addr),
    .io_chosen(rd_arb_io_chosen)
  );
  assign io_mem_aw_valid = wstate == 2'h1; // @[DME.scala 226:19]
  assign io_mem_w_valid = 1'h0; // @[DME.scala 230:18]
  assign io_mem_w_bits_last = wr_cnt == 32'h0; // @[DME.scala 232:22]
  assign io_mem_b_ready = wstate == 2'h3; // @[DME.scala 234:18]
  assign io_mem_ar_valid = rstate == 2'h1; // @[DME.scala 236:19]
  assign io_mem_ar_bits_addr = rd_addr; // @[DME.scala 237:23]
  assign io_mem_r_ready = _T_43 & _GEN_40; // @[DME.scala 240:18]
  assign io_dme_rd_0_data_valid = _T_24 & io_mem_r_valid; // @[DME.scala 215:29]
  assign io_dme_rd_0_data_bits = io_mem_r_bits_data; // @[DME.scala 216:28]
  assign io_dme_rd_1_data_valid = _T_26 & io_mem_r_valid; // @[DME.scala 215:29]
  assign io_dme_rd_1_data_bits = io_mem_r_bits_data; // @[DME.scala 216:28]
  assign io_dme_rd_2_data_valid = _T_28 & io_mem_r_valid; // @[DME.scala 215:29]
  assign io_dme_rd_2_data_bits = io_mem_r_bits_data; // @[DME.scala 216:28]
  assign rd_arb_io_in_0_valid = io_dme_rd_0_cmd_valid; // @[DME.scala 134:21]
  assign rd_arb_io_in_0_bits_addr = io_dme_rd_0_cmd_bits_addr; // @[DME.scala 134:21]
  assign rd_arb_io_in_1_valid = io_dme_rd_1_cmd_valid; // @[DME.scala 134:21]
  assign rd_arb_io_in_1_bits_addr = io_dme_rd_1_cmd_bits_addr; // @[DME.scala 134:21]
  assign rd_arb_io_in_2_valid = io_dme_rd_2_cmd_valid; // @[DME.scala 134:21]
  assign rd_arb_io_in_2_bits_addr = io_dme_rd_2_cmd_bits_addr; // @[DME.scala 134:21]
  assign rd_arb_io_out_ready = rstate == 2'h0; // @[DME.scala 210:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rd_arb_chosen = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  rstate = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  wstate = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  wr_cnt = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  rd_addr = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T) begin
      rd_arb_chosen <= rd_arb_io_chosen;
    end
    if (reset) begin
      rstate <= 2'h0;
    end else if (_T_1) begin
      if (rd_arb_io_out_valid) begin
        rstate <= 2'h1;
      end
    end else if (_T_2) begin
      if (io_mem_ar_ready) begin
        rstate <= 2'h2;
      end
    end else if (_T_3) begin
      if (_T_5) begin
        rstate <= 2'h0;
      end
    end
    if (reset) begin
      wstate <= 2'h0;
    end else if (!(_T_11)) begin
      if (_T_12) begin
        if (io_mem_aw_ready) begin
          wstate <= 2'h2;
        end
      end else if (!(_T_13)) begin
        if (_T_17) begin
          if (io_mem_b_valid) begin
            wstate <= 2'h0;
          end
        end
      end
    end
    if (reset) begin
      wr_cnt <= 32'h0;
    end else if (_T_7) begin
      wr_cnt <= 32'h0;
    end else if (_T_8) begin
      wr_cnt <= _T_10;
    end
    if (reset) begin
      rd_addr <= 32'h0;
    end else if (_T) begin
      rd_addr <= rd_arb_io_out_bits_addr;
    end
  end
endmodule
module memoryWrapper(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [7:0]  io_in_bits_inst,
  input  [63:0] io_in_bits_data,
  input  [2:0]  io_in_bits_src,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output        io_mem_b_ready,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [15:0] io_mem_ar_bits_len,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [63:0] io_out_bits_data,
  output [2:0]  io_out_bits_dst
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] addrReg; // @[mainMemWrapper.scala 36:26]
  reg [2:0] numberOfLines; // @[mainMemWrapper.scala 37:32]
  reg [2:0] srcReg; // @[mainMemWrapper.scala 38:25]
  reg [31:0] returnAddr; // @[mainMemWrapper.scala 39:29]
  reg [63:0] dataRegRead_0; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegRead_1; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegRead_2; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegRead_3; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegRead_4; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegRead_5; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegRead_6; // @[mainMemWrapper.scala 40:30]
  reg [63:0] dataRegWrite_0; // @[mainMemWrapper.scala 41:31]
  reg [2:0] stReg; // @[mainMemWrapper.scala 44:24]
  wire  _T_2 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = stReg == 3'h0; // @[mainMemWrapper.scala 47:35]
  wire  _T_4 = _T_2 & _T_3; // @[mainMemWrapper.scala 47:27]
  wire  _T_6 = io_in_bits_data[31:0] != 32'h0; // @[mainMemWrapper.scala 47:80]
  wire  start = _T_4 & _T_6; // @[mainMemWrapper.scala 47:46]
  wire [31:0] _T_9 = {io_in_bits_data[31:3], 3'h0}; // @[mainMemWrapper.scala 50:58]
  wire  _T_11 = io_in_bits_data[2:0] == 3'h0; // @[mainMemWrapper.scala 51:51]
  wire  _T_15 = io_in_bits_inst == 8'h1; // @[mainMemWrapper.scala 58:54]
  wire  writeInst = start & _T_15; // @[mainMemWrapper.scala 58:36]
  wire  _T_17 = io_mem_r_ready & io_mem_r_valid; // @[Decoupled.scala 40:37]
  reg [2:0] readCount; // @[Counter.scala 29:33]
  wire  _T_18 = readCount == 3'h6; // @[Counter.scala 38:24]
  wire [2:0] _T_20 = readCount + 3'h1; // @[Counter.scala 39:22]
  wire  writeWrapped = io_mem_w_ready & io_mem_w_valid; // @[Decoupled.scala 40:37]
  wire  _T_22 = stReg == 3'h5; // @[mainMemWrapper.scala 65:55]
  reg [19:0] dramLatencyCnt; // @[Counter.scala 29:33]
  wire  _T_24 = dramLatencyCnt == 20'hf423f; // @[Counter.scala 38:24]
  wire [19:0] _T_26 = dramLatencyCnt + 20'h1; // @[Counter.scala 39:22]
  wire  _T_27 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [19:0] nextPacket; // @[Counter.scala 29:33]
  wire  _T_29 = nextPacket == 20'hf423f; // @[Counter.scala 38:24]
  wire [19:0] _T_31 = nextPacket + 20'h1; // @[Counter.scala 39:22]
  wire [2:0] _T_33 = numberOfLines - 3'h1; // @[mainMemWrapper.scala 67:62]
  wire [19:0] _GEN_75 = {{17'd0}, _T_33}; // @[mainMemWrapper.scala 67:44]
  wire  packetsDone = nextPacket == _GEN_75; // @[mainMemWrapper.scala 67:44]
  wire [31:0] _T_38 = returnAddr + 32'h8; // @[mainMemWrapper.scala 70:34]
  wire  _T_43 = stReg == 3'h1; // @[mainMemWrapper.scala 82:38]
  wire  _T_45 = stReg == 3'h2; // @[mainMemWrapper.scala 85:37]
  wire [3:0] _T_47 = 3'h1 * numberOfLines; // @[mainMemWrapper.scala 89:35]
  wire [3:0] _T_49 = _T_47 - 4'h1; // @[mainMemWrapper.scala 89:51]
  wire [20:0] _T_51 = nextPacket * 20'h1; // @[mainMemWrapper.scala 101:78]
  wire [21:0] _T_52 = {{1'd0}, _T_51}; // @[mainMemWrapper.scala 101:88]
  wire [63:0] _GEN_34 = 3'h1 == _T_52[2:0] ? dataRegRead_1 : dataRegRead_0; // @[mainMemWrapper.scala 101:22]
  wire [63:0] _GEN_35 = 3'h2 == _T_52[2:0] ? dataRegRead_2 : _GEN_34; // @[mainMemWrapper.scala 101:22]
  wire [63:0] _GEN_36 = 3'h3 == _T_52[2:0] ? dataRegRead_3 : _GEN_35; // @[mainMemWrapper.scala 101:22]
  wire [63:0] _GEN_37 = 3'h4 == _T_52[2:0] ? dataRegRead_4 : _GEN_36; // @[mainMemWrapper.scala 101:22]
  wire [63:0] _GEN_38 = 3'h5 == _T_52[2:0] ? dataRegRead_5 : _GEN_37; // @[mainMemWrapper.scala 101:22]
  wire  _T_55 = 3'h0 == stReg; // @[Conditional.scala 37:30]
  wire  _T_56 = 3'h3 == stReg; // @[Conditional.scala 37:30]
  wire  _T_57 = io_mem_ar_ready & io_mem_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_58 = 3'h4 == stReg; // @[Conditional.scala 37:30]
  wire  _T_60 = _T_17 & io_mem_r_bits_last; // @[mainMemWrapper.scala 129:34]
  wire  _T_61 = 3'h1 == stReg; // @[Conditional.scala 37:30]
  wire  _T_62 = io_mem_aw_ready & io_mem_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_63 = 3'h2 == stReg; // @[Conditional.scala 37:30]
  wire  _T_64 = 3'h5 == stReg; // @[Conditional.scala 37:30]
  wire  _T_65 = dramLatencyCnt > 20'hc8; // @[mainMemWrapper.scala 146:34]
  wire  _T_67 = packetsDone & _T_27; // @[mainMemWrapper.scala 148:34]
  wire  _GEN_49 = _T_64 & _T_65; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_63 ? 1'h0 : _GEN_49; // @[Conditional.scala 39:67]
  wire  _GEN_56 = _T_61 ? 1'h0 : _T_63; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_61 ? 1'h0 : _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_60 = _T_58 ? 1'h0 : _T_61; // @[Conditional.scala 39:67]
  wire  _GEN_61 = _T_58 ? 1'h0 : _GEN_56; // @[Conditional.scala 39:67]
  wire  _GEN_62 = _T_58 ? 1'h0 : _GEN_57; // @[Conditional.scala 39:67]
  wire  _GEN_65 = _T_56 ? 1'h0 : _T_58; // @[Conditional.scala 39:67]
  wire  _GEN_66 = _T_56 ? 1'h0 : _GEN_60; // @[Conditional.scala 39:67]
  wire  _GEN_67 = _T_56 ? 1'h0 : _GEN_61; // @[Conditional.scala 39:67]
  wire  _GEN_68 = _T_56 ? 1'h0 : _GEN_62; // @[Conditional.scala 39:67]
  assign io_in_ready = stReg == 3'h0; // @[mainMemWrapper.scala 56:17]
  assign io_mem_aw_valid = _T_55 ? 1'h0 : _GEN_66; // @[mainMemWrapper.scala 93:21 mainMemWrapper.scala 134:29]
  assign io_mem_aw_bits_addr = _T_43 ? addrReg : 32'h0; // @[mainMemWrapper.scala 82:25]
  assign io_mem_w_valid = _T_55 ? 1'h0 : _GEN_67; // @[mainMemWrapper.scala 95:20 mainMemWrapper.scala 140:28]
  assign io_mem_w_bits_data = _T_45 ? dataRegWrite_0 : 64'h0; // @[mainMemWrapper.scala 85:24]
  assign io_mem_b_ready = stReg == 3'h2; // @[mainMemWrapper.scala 90:20]
  assign io_mem_ar_valid = _T_55 ? 1'h0 : _T_56; // @[mainMemWrapper.scala 92:21 mainMemWrapper.scala 122:29]
  assign io_mem_ar_bits_addr = addrReg; // @[mainMemWrapper.scala 88:25]
  assign io_mem_ar_bits_len = {{12'd0}, _T_49}; // @[mainMemWrapper.scala 89:24]
  assign io_mem_r_ready = _T_55 ? 1'h0 : _GEN_65; // @[mainMemWrapper.scala 94:20 mainMemWrapper.scala 128:28]
  assign io_out_valid = _T_55 ? 1'h0 : _GEN_68; // @[mainMemWrapper.scala 109:18 mainMemWrapper.scala 147:30]
  assign io_out_bits_addr = returnAddr; // @[mainMemWrapper.scala 102:22]
  assign io_out_bits_data = 3'h6 == _T_52[2:0] ? dataRegRead_6 : _GEN_38; // @[mainMemWrapper.scala 101:22]
  assign io_out_bits_dst = srcReg; // @[mainMemWrapper.scala 105:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addrReg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  numberOfLines = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  srcReg = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  returnAddr = _RAND_3[31:0];
  _RAND_4 = {2{`RANDOM}};
  dataRegRead_0 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  dataRegRead_1 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataRegRead_2 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataRegRead_3 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataRegRead_4 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  dataRegRead_5 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  dataRegRead_6 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  dataRegWrite_0 = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  stReg = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  readCount = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  dramLatencyCnt = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  nextPacket = _RAND_15[19:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addrReg <= 32'h0;
    end else if (start) begin
      addrReg <= _T_9;
    end
    if (reset) begin
      numberOfLines <= 3'h0;
    end else if (start) begin
      if (_T_11) begin
        numberOfLines <= 3'h1;
      end else begin
        numberOfLines <= io_in_bits_data[2:0];
      end
    end
    if (reset) begin
      srcReg <= 3'h0;
    end else if (start) begin
      srcReg <= io_in_bits_src;
    end
    if (reset) begin
      returnAddr <= 32'h0;
    end else if (_T_27) begin
      returnAddr <= _T_38;
    end else if (start) begin
      returnAddr <= io_in_bits_addr;
    end
    if (reset) begin
      dataRegRead_0 <= 64'h0;
    end else if (_T_17) begin
      if (3'h0 == readCount) begin
        dataRegRead_0 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegRead_1 <= 64'h0;
    end else if (_T_17) begin
      if (3'h1 == readCount) begin
        dataRegRead_1 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegRead_2 <= 64'h0;
    end else if (_T_17) begin
      if (3'h2 == readCount) begin
        dataRegRead_2 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegRead_3 <= 64'h0;
    end else if (_T_17) begin
      if (3'h3 == readCount) begin
        dataRegRead_3 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegRead_4 <= 64'h0;
    end else if (_T_17) begin
      if (3'h4 == readCount) begin
        dataRegRead_4 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegRead_5 <= 64'h0;
    end else if (_T_17) begin
      if (3'h5 == readCount) begin
        dataRegRead_5 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegRead_6 <= 64'h0;
    end else if (_T_17) begin
      if (3'h6 == readCount) begin
        dataRegRead_6 <= io_mem_r_bits_data;
      end
    end
    if (reset) begin
      dataRegWrite_0 <= 64'h0;
    end else if (writeInst) begin
      dataRegWrite_0 <= io_in_bits_data;
    end
    if (reset) begin
      stReg <= 3'h0;
    end else if (_T_55) begin
      if (start) begin
        if (writeInst) begin
          stReg <= 3'h1;
        end else begin
          stReg <= 3'h3;
        end
      end
    end else if (_T_56) begin
      if (_T_57) begin
        stReg <= 3'h4;
      end
    end else if (_T_58) begin
      if (_T_60) begin
        stReg <= 3'h5;
      end
    end else if (_T_61) begin
      if (_T_62) begin
        stReg <= 3'h2;
      end
    end else if (_T_63) begin
      if (writeWrapped) begin
        stReg <= 3'h0;
      end
    end else if (_T_64) begin
      if (_T_65) begin
        if (_T_67) begin
          stReg <= 3'h0;
        end
      end
    end
    if (reset) begin
      readCount <= 3'h0;
    end else if (start) begin
      readCount <= 3'h0;
    end else if (_T_17) begin
      if (_T_18) begin
        readCount <= 3'h0;
      end else begin
        readCount <= _T_20;
      end
    end
    if (reset) begin
      dramLatencyCnt <= 20'h0;
    end else if (start) begin
      dramLatencyCnt <= 20'h0;
    end else if (_T_22) begin
      if (_T_24) begin
        dramLatencyCnt <= 20'h0;
      end else begin
        dramLatencyCnt <= _T_26;
      end
    end
    if (reset) begin
      nextPacket <= 20'h0;
    end else if (start) begin
      nextPacket <= 20'h0;
    end else if (_T_27) begin
      if (_T_29) begin
        nextPacket <= 20'h0;
      end else begin
        nextPacket <= _T_31;
      end
    end
  end
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_inst,
  input  [63:0] io_enq_bits_data,
  input  [2:0]  io_enq_bits_src,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_inst,
  output [63:0] io_deq_bits_data,
  output [2:0]  io_deq_bits_src
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:127]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_11_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_addr__T_11_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [7:0] ram_inst [0:127]; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_11_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_inst__T_11_addr; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_3_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_inst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:127]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_11_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_data__T_11_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_src [0:127]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_src__T_11_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_src__T_11_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_src__T_3_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_src__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_en; // @[Decoupled.scala 209:16]
  reg [6:0] enq_ptr_value; // @[Counter.scala 29:33]
  reg [6:0] deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [6:0] _T_5 = enq_ptr_value + 7'h1; // @[Counter.scala 39:22]
  wire [6:0] _T_7 = deq_ptr_value + 7'h1; // @[Counter.scala 39:22]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram_addr__T_11_addr = deq_ptr_value;
  assign ram_addr__T_11_data = ram_addr[ram_addr__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_3_data = io_enq_bits_addr;
  assign ram_addr__T_3_addr = enq_ptr_value;
  assign ram_addr__T_3_mask = 1'h1;
  assign ram_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst__T_11_addr = deq_ptr_value;
  assign ram_inst__T_11_data = ram_inst[ram_inst__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst__T_3_data = io_enq_bits_inst;
  assign ram_inst__T_3_addr = enq_ptr_value;
  assign ram_inst__T_3_mask = 1'h1;
  assign ram_inst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_11_addr = deq_ptr_value;
  assign ram_data__T_11_data = ram_data[ram_data__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = enq_ptr_value;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_src__T_11_addr = deq_ptr_value;
  assign ram_src__T_11_data = ram_src[ram_src__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_src__T_3_data = io_enq_bits_src;
  assign ram_src__T_3_addr = enq_ptr_value;
  assign ram_src__T_3_mask = 1'h1;
  assign ram_src__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst = ram_inst__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_src = ram_src__T_11_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_inst[initvar] = _RAND_1[7:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_src[initvar] = _RAND_3[2:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enq_ptr_value = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  deq_ptr_value = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  maybe_full = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_3_en & ram_addr__T_3_mask) begin
      ram_addr[ram_addr__T_3_addr] <= ram_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst__T_3_en & ram_inst__T_3_mask) begin
      ram_inst[ram_inst__T_3_addr] <= ram_inst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_src__T_3_en & ram_src__T_3_mask) begin
      ram_src[ram_src__T_3_addr] <= ram_src__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 7'h0;
    end else if (do_enq) begin
      enq_ptr_value <= _T_5;
    end
    if (reset) begin
      deq_ptr_value <= 7'h0;
    end else if (do_deq) begin
      deq_ptr_value <= _T_7;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_inst,
  input  [63:0] io_enq_bits_data,
  input  [2:0]  io_enq_bits_src,
  input  [2:0]  io_enq_bits_dst,
  input  [1:0]  io_enq_bits_msgType,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_inst,
  output [63:0] io_deq_bits_data,
  output [2:0]  io_deq_bits_src,
  output [2:0]  io_deq_bits_dst,
  output [1:0]  io_deq_bits_msgType
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:1]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_11_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [7:0] ram_inst [0:1]; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_11_addr; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_11_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_src [0:1]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_src__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_src__T_11_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_src__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_dst [0:1]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_dst__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_11_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_dst__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_3_en; // @[Decoupled.scala 209:16]
  reg [1:0] ram_msgType [0:1]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_msgType__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_11_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_msgType__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_3_en; // @[Decoupled.scala 209:16]
  reg  enq_ptr_value; // @[Counter.scala 29:33]
  reg  deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = enq_ptr_value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_7 = deq_ptr_value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  wire  _T_10 = ~full; // @[Decoupled.scala 232:19]
  assign ram_addr__T_11_addr = deq_ptr_value;
  assign ram_addr__T_11_data = ram_addr[ram_addr__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_3_data = io_enq_bits_addr;
  assign ram_addr__T_3_addr = enq_ptr_value;
  assign ram_addr__T_3_mask = 1'h1;
  assign ram_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst__T_11_addr = deq_ptr_value;
  assign ram_inst__T_11_data = ram_inst[ram_inst__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst__T_3_data = io_enq_bits_inst;
  assign ram_inst__T_3_addr = enq_ptr_value;
  assign ram_inst__T_3_mask = 1'h1;
  assign ram_inst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_11_addr = deq_ptr_value;
  assign ram_data__T_11_data = ram_data[ram_data__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = enq_ptr_value;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_src__T_11_addr = deq_ptr_value;
  assign ram_src__T_11_data = ram_src[ram_src__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_src__T_3_data = io_enq_bits_src;
  assign ram_src__T_3_addr = enq_ptr_value;
  assign ram_src__T_3_mask = 1'h1;
  assign ram_src__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_dst__T_11_addr = deq_ptr_value;
  assign ram_dst__T_11_data = ram_dst[ram_dst__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_dst__T_3_data = io_enq_bits_dst;
  assign ram_dst__T_3_addr = enq_ptr_value;
  assign ram_dst__T_3_mask = 1'h1;
  assign ram_dst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_msgType__T_11_addr = deq_ptr_value;
  assign ram_msgType__T_11_data = ram_msgType[ram_msgType__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_msgType__T_3_data = io_enq_bits_msgType;
  assign ram_msgType__T_3_addr = enq_ptr_value;
  assign ram_msgType__T_3_mask = 1'h1;
  assign ram_msgType__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | _T_10; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst = ram_inst__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_src = ram_src__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_dst = ram_dst__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_msgType = ram_msgType__T_11_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_inst[initvar] = _RAND_1[7:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_src[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_dst[initvar] = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_msgType[initvar] = _RAND_5[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enq_ptr_value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  deq_ptr_value = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_3_en & ram_addr__T_3_mask) begin
      ram_addr[ram_addr__T_3_addr] <= ram_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst__T_3_en & ram_inst__T_3_mask) begin
      ram_inst[ram_inst__T_3_addr] <= ram_inst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_src__T_3_en & ram_src__T_3_mask) begin
      ram_src[ram_src__T_3_addr] <= ram_src__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_dst__T_3_en & ram_dst__T_3_mask) begin
      ram_dst[ram_dst__T_3_addr] <= ram_dst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_msgType__T_3_en & ram_msgType__T_3_mask) begin
      ram_msgType[ram_msgType__T_3_addr] <= ram_msgType__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 1'h0;
    end else if (do_enq) begin
      enq_ptr_value <= _T_5;
    end
    if (reset) begin
      deq_ptr_value <= 1'h0;
    end else if (do_deq) begin
      deq_ptr_value <= _T_7;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_3(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_inst,
  input  [63:0] io_enq_bits_data,
  input  [2:0]  io_enq_bits_src,
  input  [2:0]  io_enq_bits_dst,
  input  [1:0]  io_enq_bits_msgType,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_inst,
  output [63:0] io_deq_bits_data,
  output [2:0]  io_deq_bits_src,
  output [2:0]  io_deq_bits_dst,
  output [1:0]  io_deq_bits_msgType
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:1]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_11_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [7:0] ram_inst [0:1]; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_11_addr; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_11_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_src [0:1]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_src__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_src__T_11_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_src__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_src__T_3_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_dst [0:1]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_dst__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_11_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_dst__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_dst__T_3_en; // @[Decoupled.scala 209:16]
  reg [1:0] ram_msgType [0:1]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_msgType__T_11_data; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_11_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_msgType__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_msgType__T_3_en; // @[Decoupled.scala 209:16]
  reg  enq_ptr_value; // @[Counter.scala 29:33]
  reg  deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = enq_ptr_value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_7 = deq_ptr_value + 1'h1; // @[Counter.scala 39:22]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram_addr__T_11_addr = deq_ptr_value;
  assign ram_addr__T_11_data = ram_addr[ram_addr__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_3_data = io_enq_bits_addr;
  assign ram_addr__T_3_addr = enq_ptr_value;
  assign ram_addr__T_3_mask = 1'h1;
  assign ram_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst__T_11_addr = deq_ptr_value;
  assign ram_inst__T_11_data = ram_inst[ram_inst__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst__T_3_data = io_enq_bits_inst;
  assign ram_inst__T_3_addr = enq_ptr_value;
  assign ram_inst__T_3_mask = 1'h1;
  assign ram_inst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_11_addr = deq_ptr_value;
  assign ram_data__T_11_data = ram_data[ram_data__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = enq_ptr_value;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_src__T_11_addr = deq_ptr_value;
  assign ram_src__T_11_data = ram_src[ram_src__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_src__T_3_data = io_enq_bits_src;
  assign ram_src__T_3_addr = enq_ptr_value;
  assign ram_src__T_3_mask = 1'h1;
  assign ram_src__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_dst__T_11_addr = deq_ptr_value;
  assign ram_dst__T_11_data = ram_dst[ram_dst__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_dst__T_3_data = io_enq_bits_dst;
  assign ram_dst__T_3_addr = enq_ptr_value;
  assign ram_dst__T_3_mask = 1'h1;
  assign ram_dst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_msgType__T_11_addr = deq_ptr_value;
  assign ram_msgType__T_11_data = ram_msgType[ram_msgType__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_msgType__T_3_data = io_enq_bits_msgType;
  assign ram_msgType__T_3_addr = enq_ptr_value;
  assign ram_msgType__T_3_mask = 1'h1;
  assign ram_msgType__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst = ram_inst__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_src = ram_src__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_dst = ram_dst__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_msgType = ram_msgType__T_11_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_inst[initvar] = _RAND_1[7:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_src[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_dst[initvar] = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_msgType[initvar] = _RAND_5[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enq_ptr_value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  deq_ptr_value = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_3_en & ram_addr__T_3_mask) begin
      ram_addr[ram_addr__T_3_addr] <= ram_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst__T_3_en & ram_inst__T_3_mask) begin
      ram_inst[ram_inst__T_3_addr] <= ram_inst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_src__T_3_en & ram_src__T_3_mask) begin
      ram_src[ram_src__T_3_addr] <= ram_src__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_dst__T_3_en & ram_dst__T_3_mask) begin
      ram_dst[ram_dst__T_3_addr] <= ram_dst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_msgType__T_3_en & ram_msgType__T_3_mask) begin
      ram_msgType[ram_msgType__T_3_addr] <= ram_msgType__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 1'h0;
    end else if (do_enq) begin
      enq_ptr_value <= _T_5;
    end
    if (reset) begin
      deq_ptr_value <= 1'h0;
    end else if (do_deq) begin
      deq_ptr_value <= _T_7;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module RRArbiter(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [7:0]  io_in_0_bits_inst,
  input  [63:0] io_in_0_bits_data,
  input  [2:0]  io_in_0_bits_src,
  input  [2:0]  io_in_0_bits_dst,
  input  [1:0]  io_in_0_bits_msgType,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [7:0]  io_in_1_bits_inst,
  input  [63:0] io_in_1_bits_data,
  input  [2:0]  io_in_1_bits_src,
  input  [2:0]  io_in_1_bits_dst,
  input  [1:0]  io_in_1_bits_msgType,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [7:0]  io_out_bits_inst,
  output [63:0] io_out_bits_data,
  output [2:0]  io_out_bits_src,
  output [2:0]  io_out_bits_dst,
  output [1:0]  io_out_bits_msgType,
  output        io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  lastGrant; // @[Reg.scala 15:16]
  wire  grantMask_1 = 1'h1 > lastGrant; // @[Arbiter.scala 67:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbiter.scala 68:75]
  wire  _T_2 = validMask_1 | io_in_0_valid; // @[Arbiter.scala 31:68]
  wire  _T_4 = ~validMask_1; // @[Arbiter.scala 31:78]
  wire  _T_5 = ~_T_2; // @[Arbiter.scala 31:78]
  wire  _T_9 = grantMask_1 | _T_5; // @[Arbiter.scala 72:50]
  wire  _GEN_17 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_4 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_9 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:15]
  assign io_out_bits_inst = io_chosen ? io_in_1_bits_inst : io_in_0_bits_inst; // @[Arbiter.scala 42:15]
  assign io_out_bits_data = io_chosen ? io_in_1_bits_data : io_in_0_bits_data; // @[Arbiter.scala 42:15]
  assign io_out_bits_src = io_chosen ? io_in_1_bits_src : io_in_0_bits_src; // @[Arbiter.scala 42:15]
  assign io_out_bits_dst = io_chosen ? io_in_1_bits_dst : io_in_0_bits_dst; // @[Arbiter.scala 42:15]
  assign io_out_bits_msgType = io_chosen ? io_in_1_bits_msgType : io_in_0_bits_msgType; // @[Arbiter.scala 42:15]
  assign io_chosen = validMask_1 | _GEN_17; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T) begin
      lastGrant <= io_chosen;
    end
  end
endmodule
module Router(
  input         clock,
  input         reset,
  input         io_cacheIn_valid,
  input  [31:0] io_cacheIn_bits_addr,
  input  [7:0]  io_cacheIn_bits_inst,
  input  [63:0] io_cacheIn_bits_data,
  input         io_cacheOut_ready,
  output        io_cacheOut_valid,
  output [31:0] io_cacheOut_bits_addr,
  output [7:0]  io_cacheOut_bits_inst,
  output [63:0] io_cacheOut_bits_data,
  output [1:0]  io_cacheOut_bits_msgType,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [7:0]  io_in_bits_inst,
  input  [63:0] io_in_bits_data,
  input  [2:0]  io_in_bits_src,
  input  [2:0]  io_in_bits_dst,
  input  [1:0]  io_in_bits_msgType,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [7:0]  io_out_bits_inst,
  output [63:0] io_out_bits_data,
  output [2:0]  io_out_bits_src,
  output [2:0]  io_out_bits_dst,
  output [1:0]  io_out_bits_msgType
);
  wire  cache_in_Q_clock; // @[Router.scala 19:26]
  wire  cache_in_Q_reset; // @[Router.scala 19:26]
  wire  cache_in_Q_io_enq_ready; // @[Router.scala 19:26]
  wire  cache_in_Q_io_enq_valid; // @[Router.scala 19:26]
  wire [31:0] cache_in_Q_io_enq_bits_addr; // @[Router.scala 19:26]
  wire [7:0] cache_in_Q_io_enq_bits_inst; // @[Router.scala 19:26]
  wire [63:0] cache_in_Q_io_enq_bits_data; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_enq_bits_src; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_enq_bits_dst; // @[Router.scala 19:26]
  wire [1:0] cache_in_Q_io_enq_bits_msgType; // @[Router.scala 19:26]
  wire  cache_in_Q_io_deq_ready; // @[Router.scala 19:26]
  wire  cache_in_Q_io_deq_valid; // @[Router.scala 19:26]
  wire [31:0] cache_in_Q_io_deq_bits_addr; // @[Router.scala 19:26]
  wire [7:0] cache_in_Q_io_deq_bits_inst; // @[Router.scala 19:26]
  wire [63:0] cache_in_Q_io_deq_bits_data; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_deq_bits_src; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_deq_bits_dst; // @[Router.scala 19:26]
  wire [1:0] cache_in_Q_io_deq_bits_msgType; // @[Router.scala 19:26]
  wire  cache_out_Q_clock; // @[Router.scala 20:27]
  wire  cache_out_Q_reset; // @[Router.scala 20:27]
  wire  cache_out_Q_io_enq_ready; // @[Router.scala 20:27]
  wire  cache_out_Q_io_enq_valid; // @[Router.scala 20:27]
  wire [31:0] cache_out_Q_io_enq_bits_addr; // @[Router.scala 20:27]
  wire [7:0] cache_out_Q_io_enq_bits_inst; // @[Router.scala 20:27]
  wire [63:0] cache_out_Q_io_enq_bits_data; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_enq_bits_src; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_enq_bits_dst; // @[Router.scala 20:27]
  wire [1:0] cache_out_Q_io_enq_bits_msgType; // @[Router.scala 20:27]
  wire  cache_out_Q_io_deq_ready; // @[Router.scala 20:27]
  wire  cache_out_Q_io_deq_valid; // @[Router.scala 20:27]
  wire [31:0] cache_out_Q_io_deq_bits_addr; // @[Router.scala 20:27]
  wire [7:0] cache_out_Q_io_deq_bits_inst; // @[Router.scala 20:27]
  wire [63:0] cache_out_Q_io_deq_bits_data; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_deq_bits_src; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_deq_bits_dst; // @[Router.scala 20:27]
  wire [1:0] cache_out_Q_io_deq_bits_msgType; // @[Router.scala 20:27]
  wire  in_Q_clock; // @[Router.scala 21:20]
  wire  in_Q_reset; // @[Router.scala 21:20]
  wire  in_Q_io_enq_ready; // @[Router.scala 21:20]
  wire  in_Q_io_enq_valid; // @[Router.scala 21:20]
  wire [31:0] in_Q_io_enq_bits_addr; // @[Router.scala 21:20]
  wire [7:0] in_Q_io_enq_bits_inst; // @[Router.scala 21:20]
  wire [63:0] in_Q_io_enq_bits_data; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_enq_bits_src; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_enq_bits_dst; // @[Router.scala 21:20]
  wire [1:0] in_Q_io_enq_bits_msgType; // @[Router.scala 21:20]
  wire  in_Q_io_deq_ready; // @[Router.scala 21:20]
  wire  in_Q_io_deq_valid; // @[Router.scala 21:20]
  wire [31:0] in_Q_io_deq_bits_addr; // @[Router.scala 21:20]
  wire [7:0] in_Q_io_deq_bits_inst; // @[Router.scala 21:20]
  wire [63:0] in_Q_io_deq_bits_data; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_deq_bits_src; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_deq_bits_dst; // @[Router.scala 21:20]
  wire [1:0] in_Q_io_deq_bits_msgType; // @[Router.scala 21:20]
  wire  arbiter_clock; // @[Router.scala 23:23]
  wire  arbiter_io_in_0_ready; // @[Router.scala 23:23]
  wire  arbiter_io_in_0_valid; // @[Router.scala 23:23]
  wire [31:0] arbiter_io_in_0_bits_addr; // @[Router.scala 23:23]
  wire [7:0] arbiter_io_in_0_bits_inst; // @[Router.scala 23:23]
  wire [63:0] arbiter_io_in_0_bits_data; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_0_bits_src; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_0_bits_dst; // @[Router.scala 23:23]
  wire [1:0] arbiter_io_in_0_bits_msgType; // @[Router.scala 23:23]
  wire  arbiter_io_in_1_ready; // @[Router.scala 23:23]
  wire  arbiter_io_in_1_valid; // @[Router.scala 23:23]
  wire [31:0] arbiter_io_in_1_bits_addr; // @[Router.scala 23:23]
  wire [7:0] arbiter_io_in_1_bits_inst; // @[Router.scala 23:23]
  wire [63:0] arbiter_io_in_1_bits_data; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_1_bits_src; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_1_bits_dst; // @[Router.scala 23:23]
  wire [1:0] arbiter_io_in_1_bits_msgType; // @[Router.scala 23:23]
  wire  arbiter_io_out_ready; // @[Router.scala 23:23]
  wire  arbiter_io_out_valid; // @[Router.scala 23:23]
  wire [31:0] arbiter_io_out_bits_addr; // @[Router.scala 23:23]
  wire [7:0] arbiter_io_out_bits_inst; // @[Router.scala 23:23]
  wire [63:0] arbiter_io_out_bits_data; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_out_bits_src; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_out_bits_dst; // @[Router.scala 23:23]
  wire [1:0] arbiter_io_out_bits_msgType; // @[Router.scala 23:23]
  wire  arbiter_io_chosen; // @[Router.scala 23:23]
  wire  _T = in_Q_io_deq_bits_dst == 3'h0; // @[Router.scala 34:74]
  wire  _T_2 = in_Q_io_deq_bits_dst != 3'h0; // @[Router.scala 37:72]
  wire  _T_5 = arbiter_io_in_1_ready & _T_2; // @[Router.scala 38:48]
  wire  _T_7 = cache_out_Q_io_enq_ready & _T; // @[Router.scala 38:113]
  Queue_1 cache_in_Q ( // @[Router.scala 19:26]
    .clock(cache_in_Q_clock),
    .reset(cache_in_Q_reset),
    .io_enq_ready(cache_in_Q_io_enq_ready),
    .io_enq_valid(cache_in_Q_io_enq_valid),
    .io_enq_bits_addr(cache_in_Q_io_enq_bits_addr),
    .io_enq_bits_inst(cache_in_Q_io_enq_bits_inst),
    .io_enq_bits_data(cache_in_Q_io_enq_bits_data),
    .io_enq_bits_src(cache_in_Q_io_enq_bits_src),
    .io_enq_bits_dst(cache_in_Q_io_enq_bits_dst),
    .io_enq_bits_msgType(cache_in_Q_io_enq_bits_msgType),
    .io_deq_ready(cache_in_Q_io_deq_ready),
    .io_deq_valid(cache_in_Q_io_deq_valid),
    .io_deq_bits_addr(cache_in_Q_io_deq_bits_addr),
    .io_deq_bits_inst(cache_in_Q_io_deq_bits_inst),
    .io_deq_bits_data(cache_in_Q_io_deq_bits_data),
    .io_deq_bits_src(cache_in_Q_io_deq_bits_src),
    .io_deq_bits_dst(cache_in_Q_io_deq_bits_dst),
    .io_deq_bits_msgType(cache_in_Q_io_deq_bits_msgType)
  );
  Queue_1 cache_out_Q ( // @[Router.scala 20:27]
    .clock(cache_out_Q_clock),
    .reset(cache_out_Q_reset),
    .io_enq_ready(cache_out_Q_io_enq_ready),
    .io_enq_valid(cache_out_Q_io_enq_valid),
    .io_enq_bits_addr(cache_out_Q_io_enq_bits_addr),
    .io_enq_bits_inst(cache_out_Q_io_enq_bits_inst),
    .io_enq_bits_data(cache_out_Q_io_enq_bits_data),
    .io_enq_bits_src(cache_out_Q_io_enq_bits_src),
    .io_enq_bits_dst(cache_out_Q_io_enq_bits_dst),
    .io_enq_bits_msgType(cache_out_Q_io_enq_bits_msgType),
    .io_deq_ready(cache_out_Q_io_deq_ready),
    .io_deq_valid(cache_out_Q_io_deq_valid),
    .io_deq_bits_addr(cache_out_Q_io_deq_bits_addr),
    .io_deq_bits_inst(cache_out_Q_io_deq_bits_inst),
    .io_deq_bits_data(cache_out_Q_io_deq_bits_data),
    .io_deq_bits_src(cache_out_Q_io_deq_bits_src),
    .io_deq_bits_dst(cache_out_Q_io_deq_bits_dst),
    .io_deq_bits_msgType(cache_out_Q_io_deq_bits_msgType)
  );
  Queue_3 in_Q ( // @[Router.scala 21:20]
    .clock(in_Q_clock),
    .reset(in_Q_reset),
    .io_enq_ready(in_Q_io_enq_ready),
    .io_enq_valid(in_Q_io_enq_valid),
    .io_enq_bits_addr(in_Q_io_enq_bits_addr),
    .io_enq_bits_inst(in_Q_io_enq_bits_inst),
    .io_enq_bits_data(in_Q_io_enq_bits_data),
    .io_enq_bits_src(in_Q_io_enq_bits_src),
    .io_enq_bits_dst(in_Q_io_enq_bits_dst),
    .io_enq_bits_msgType(in_Q_io_enq_bits_msgType),
    .io_deq_ready(in_Q_io_deq_ready),
    .io_deq_valid(in_Q_io_deq_valid),
    .io_deq_bits_addr(in_Q_io_deq_bits_addr),
    .io_deq_bits_inst(in_Q_io_deq_bits_inst),
    .io_deq_bits_data(in_Q_io_deq_bits_data),
    .io_deq_bits_src(in_Q_io_deq_bits_src),
    .io_deq_bits_dst(in_Q_io_deq_bits_dst),
    .io_deq_bits_msgType(in_Q_io_deq_bits_msgType)
  );
  RRArbiter arbiter ( // @[Router.scala 23:23]
    .clock(arbiter_clock),
    .io_in_0_ready(arbiter_io_in_0_ready),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_addr(arbiter_io_in_0_bits_addr),
    .io_in_0_bits_inst(arbiter_io_in_0_bits_inst),
    .io_in_0_bits_data(arbiter_io_in_0_bits_data),
    .io_in_0_bits_src(arbiter_io_in_0_bits_src),
    .io_in_0_bits_dst(arbiter_io_in_0_bits_dst),
    .io_in_0_bits_msgType(arbiter_io_in_0_bits_msgType),
    .io_in_1_ready(arbiter_io_in_1_ready),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_addr(arbiter_io_in_1_bits_addr),
    .io_in_1_bits_inst(arbiter_io_in_1_bits_inst),
    .io_in_1_bits_data(arbiter_io_in_1_bits_data),
    .io_in_1_bits_src(arbiter_io_in_1_bits_src),
    .io_in_1_bits_dst(arbiter_io_in_1_bits_dst),
    .io_in_1_bits_msgType(arbiter_io_in_1_bits_msgType),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_addr(arbiter_io_out_bits_addr),
    .io_out_bits_inst(arbiter_io_out_bits_inst),
    .io_out_bits_data(arbiter_io_out_bits_data),
    .io_out_bits_src(arbiter_io_out_bits_src),
    .io_out_bits_dst(arbiter_io_out_bits_dst),
    .io_out_bits_msgType(arbiter_io_out_bits_msgType),
    .io_chosen(arbiter_io_chosen)
  );
  assign io_cacheOut_valid = cache_out_Q_io_deq_valid; // @[Router.scala 26:15]
  assign io_cacheOut_bits_addr = cache_out_Q_io_deq_bits_addr; // @[Router.scala 26:15]
  assign io_cacheOut_bits_inst = cache_out_Q_io_deq_bits_inst; // @[Router.scala 26:15]
  assign io_cacheOut_bits_data = cache_out_Q_io_deq_bits_data; // @[Router.scala 26:15]
  assign io_cacheOut_bits_msgType = cache_out_Q_io_deq_bits_msgType; // @[Router.scala 26:15]
  assign io_in_ready = in_Q_io_enq_ready; // @[Router.scala 27:15]
  assign io_out_valid = arbiter_io_out_valid; // @[Router.scala 29:10]
  assign io_out_bits_addr = arbiter_io_out_bits_addr; // @[Router.scala 29:10]
  assign io_out_bits_inst = arbiter_io_out_bits_inst; // @[Router.scala 29:10]
  assign io_out_bits_data = arbiter_io_out_bits_data; // @[Router.scala 29:10]
  assign io_out_bits_src = arbiter_io_out_bits_src; // @[Router.scala 29:10]
  assign io_out_bits_dst = arbiter_io_out_bits_dst; // @[Router.scala 29:10]
  assign io_out_bits_msgType = arbiter_io_out_bits_msgType; // @[Router.scala 29:10]
  assign cache_in_Q_clock = clock;
  assign cache_in_Q_reset = reset;
  assign cache_in_Q_io_enq_valid = io_cacheIn_valid; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_addr = io_cacheIn_bits_addr; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_inst = io_cacheIn_bits_inst; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_data = io_cacheIn_bits_data; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_src = 3'h0; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_dst = 3'h1; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_msgType = 2'h0; // @[Router.scala 25:21]
  assign cache_in_Q_io_deq_ready = arbiter_io_in_0_ready; // @[Router.scala 31:20]
  assign cache_out_Q_clock = clock;
  assign cache_out_Q_reset = reset;
  assign cache_out_Q_io_enq_valid = in_Q_io_deq_valid & _T; // @[Router.scala 34:28]
  assign cache_out_Q_io_enq_bits_addr = in_Q_io_deq_bits_addr; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_inst = in_Q_io_deq_bits_inst; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_data = in_Q_io_deq_bits_data; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_src = in_Q_io_deq_bits_src; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_dst = in_Q_io_deq_bits_dst; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_msgType = in_Q_io_deq_bits_msgType; // @[Router.scala 33:27]
  assign cache_out_Q_io_deq_ready = io_cacheOut_ready; // @[Router.scala 26:15]
  assign in_Q_clock = clock;
  assign in_Q_reset = reset;
  assign in_Q_io_enq_valid = io_in_valid; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_addr = io_in_bits_addr; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_inst = io_in_bits_inst; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_data = io_in_bits_data; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_src = io_in_bits_src; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_dst = io_in_bits_dst; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_msgType = io_in_bits_msgType; // @[Router.scala 27:15]
  assign in_Q_io_deq_ready = _T_5 | _T_7; // @[Router.scala 38:21]
  assign arbiter_clock = clock;
  assign arbiter_io_in_0_valid = cache_in_Q_io_deq_valid; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_addr = cache_in_Q_io_deq_bits_addr; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_inst = cache_in_Q_io_deq_bits_inst; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_data = cache_in_Q_io_deq_bits_data; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_src = cache_in_Q_io_deq_bits_src; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_dst = cache_in_Q_io_deq_bits_dst; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_msgType = cache_in_Q_io_deq_bits_msgType; // @[Router.scala 31:20]
  assign arbiter_io_in_1_valid = in_Q_io_deq_valid & _T_2; // @[Router.scala 37:26]
  assign arbiter_io_in_1_bits_addr = in_Q_io_deq_bits_addr; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_inst = in_Q_io_deq_bits_inst; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_data = in_Q_io_deq_bits_data; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_src = in_Q_io_deq_bits_src; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_dst = in_Q_io_deq_bits_dst; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_msgType = in_Q_io_deq_bits_msgType; // @[Router.scala 36:25]
  assign arbiter_io_out_ready = io_out_ready; // @[Router.scala 29:10]
endmodule
module Router_1(
  input         clock,
  input         reset,
  output        io_cacheIn_ready,
  input         io_cacheIn_valid,
  input  [31:0] io_cacheIn_bits_addr,
  input  [63:0] io_cacheIn_bits_data,
  input  [2:0]  io_cacheIn_bits_dst,
  input         io_cacheOut_ready,
  output        io_cacheOut_valid,
  output [31:0] io_cacheOut_bits_addr,
  output [7:0]  io_cacheOut_bits_inst,
  output [63:0] io_cacheOut_bits_data,
  output [2:0]  io_cacheOut_bits_src,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [7:0]  io_in_bits_inst,
  input  [63:0] io_in_bits_data,
  input  [2:0]  io_in_bits_src,
  input  [2:0]  io_in_bits_dst,
  input  [1:0]  io_in_bits_msgType,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [7:0]  io_out_bits_inst,
  output [63:0] io_out_bits_data,
  output [2:0]  io_out_bits_src,
  output [2:0]  io_out_bits_dst,
  output [1:0]  io_out_bits_msgType
);
  wire  cache_in_Q_clock; // @[Router.scala 19:26]
  wire  cache_in_Q_reset; // @[Router.scala 19:26]
  wire  cache_in_Q_io_enq_ready; // @[Router.scala 19:26]
  wire  cache_in_Q_io_enq_valid; // @[Router.scala 19:26]
  wire [31:0] cache_in_Q_io_enq_bits_addr; // @[Router.scala 19:26]
  wire [7:0] cache_in_Q_io_enq_bits_inst; // @[Router.scala 19:26]
  wire [63:0] cache_in_Q_io_enq_bits_data; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_enq_bits_src; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_enq_bits_dst; // @[Router.scala 19:26]
  wire [1:0] cache_in_Q_io_enq_bits_msgType; // @[Router.scala 19:26]
  wire  cache_in_Q_io_deq_ready; // @[Router.scala 19:26]
  wire  cache_in_Q_io_deq_valid; // @[Router.scala 19:26]
  wire [31:0] cache_in_Q_io_deq_bits_addr; // @[Router.scala 19:26]
  wire [7:0] cache_in_Q_io_deq_bits_inst; // @[Router.scala 19:26]
  wire [63:0] cache_in_Q_io_deq_bits_data; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_deq_bits_src; // @[Router.scala 19:26]
  wire [2:0] cache_in_Q_io_deq_bits_dst; // @[Router.scala 19:26]
  wire [1:0] cache_in_Q_io_deq_bits_msgType; // @[Router.scala 19:26]
  wire  cache_out_Q_clock; // @[Router.scala 20:27]
  wire  cache_out_Q_reset; // @[Router.scala 20:27]
  wire  cache_out_Q_io_enq_ready; // @[Router.scala 20:27]
  wire  cache_out_Q_io_enq_valid; // @[Router.scala 20:27]
  wire [31:0] cache_out_Q_io_enq_bits_addr; // @[Router.scala 20:27]
  wire [7:0] cache_out_Q_io_enq_bits_inst; // @[Router.scala 20:27]
  wire [63:0] cache_out_Q_io_enq_bits_data; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_enq_bits_src; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_enq_bits_dst; // @[Router.scala 20:27]
  wire [1:0] cache_out_Q_io_enq_bits_msgType; // @[Router.scala 20:27]
  wire  cache_out_Q_io_deq_ready; // @[Router.scala 20:27]
  wire  cache_out_Q_io_deq_valid; // @[Router.scala 20:27]
  wire [31:0] cache_out_Q_io_deq_bits_addr; // @[Router.scala 20:27]
  wire [7:0] cache_out_Q_io_deq_bits_inst; // @[Router.scala 20:27]
  wire [63:0] cache_out_Q_io_deq_bits_data; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_deq_bits_src; // @[Router.scala 20:27]
  wire [2:0] cache_out_Q_io_deq_bits_dst; // @[Router.scala 20:27]
  wire [1:0] cache_out_Q_io_deq_bits_msgType; // @[Router.scala 20:27]
  wire  in_Q_clock; // @[Router.scala 21:20]
  wire  in_Q_reset; // @[Router.scala 21:20]
  wire  in_Q_io_enq_ready; // @[Router.scala 21:20]
  wire  in_Q_io_enq_valid; // @[Router.scala 21:20]
  wire [31:0] in_Q_io_enq_bits_addr; // @[Router.scala 21:20]
  wire [7:0] in_Q_io_enq_bits_inst; // @[Router.scala 21:20]
  wire [63:0] in_Q_io_enq_bits_data; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_enq_bits_src; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_enq_bits_dst; // @[Router.scala 21:20]
  wire [1:0] in_Q_io_enq_bits_msgType; // @[Router.scala 21:20]
  wire  in_Q_io_deq_ready; // @[Router.scala 21:20]
  wire  in_Q_io_deq_valid; // @[Router.scala 21:20]
  wire [31:0] in_Q_io_deq_bits_addr; // @[Router.scala 21:20]
  wire [7:0] in_Q_io_deq_bits_inst; // @[Router.scala 21:20]
  wire [63:0] in_Q_io_deq_bits_data; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_deq_bits_src; // @[Router.scala 21:20]
  wire [2:0] in_Q_io_deq_bits_dst; // @[Router.scala 21:20]
  wire [1:0] in_Q_io_deq_bits_msgType; // @[Router.scala 21:20]
  wire  arbiter_clock; // @[Router.scala 23:23]
  wire  arbiter_io_in_0_ready; // @[Router.scala 23:23]
  wire  arbiter_io_in_0_valid; // @[Router.scala 23:23]
  wire [31:0] arbiter_io_in_0_bits_addr; // @[Router.scala 23:23]
  wire [7:0] arbiter_io_in_0_bits_inst; // @[Router.scala 23:23]
  wire [63:0] arbiter_io_in_0_bits_data; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_0_bits_src; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_0_bits_dst; // @[Router.scala 23:23]
  wire [1:0] arbiter_io_in_0_bits_msgType; // @[Router.scala 23:23]
  wire  arbiter_io_in_1_ready; // @[Router.scala 23:23]
  wire  arbiter_io_in_1_valid; // @[Router.scala 23:23]
  wire [31:0] arbiter_io_in_1_bits_addr; // @[Router.scala 23:23]
  wire [7:0] arbiter_io_in_1_bits_inst; // @[Router.scala 23:23]
  wire [63:0] arbiter_io_in_1_bits_data; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_1_bits_src; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_in_1_bits_dst; // @[Router.scala 23:23]
  wire [1:0] arbiter_io_in_1_bits_msgType; // @[Router.scala 23:23]
  wire  arbiter_io_out_ready; // @[Router.scala 23:23]
  wire  arbiter_io_out_valid; // @[Router.scala 23:23]
  wire [31:0] arbiter_io_out_bits_addr; // @[Router.scala 23:23]
  wire [7:0] arbiter_io_out_bits_inst; // @[Router.scala 23:23]
  wire [63:0] arbiter_io_out_bits_data; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_out_bits_src; // @[Router.scala 23:23]
  wire [2:0] arbiter_io_out_bits_dst; // @[Router.scala 23:23]
  wire [1:0] arbiter_io_out_bits_msgType; // @[Router.scala 23:23]
  wire  arbiter_io_chosen; // @[Router.scala 23:23]
  wire  _T = in_Q_io_deq_bits_dst == 3'h1; // @[Router.scala 34:74]
  wire  _T_2 = in_Q_io_deq_bits_dst != 3'h1; // @[Router.scala 37:72]
  wire  _T_5 = arbiter_io_in_1_ready & _T_2; // @[Router.scala 38:48]
  wire  _T_7 = cache_out_Q_io_enq_ready & _T; // @[Router.scala 38:113]
  Queue_1 cache_in_Q ( // @[Router.scala 19:26]
    .clock(cache_in_Q_clock),
    .reset(cache_in_Q_reset),
    .io_enq_ready(cache_in_Q_io_enq_ready),
    .io_enq_valid(cache_in_Q_io_enq_valid),
    .io_enq_bits_addr(cache_in_Q_io_enq_bits_addr),
    .io_enq_bits_inst(cache_in_Q_io_enq_bits_inst),
    .io_enq_bits_data(cache_in_Q_io_enq_bits_data),
    .io_enq_bits_src(cache_in_Q_io_enq_bits_src),
    .io_enq_bits_dst(cache_in_Q_io_enq_bits_dst),
    .io_enq_bits_msgType(cache_in_Q_io_enq_bits_msgType),
    .io_deq_ready(cache_in_Q_io_deq_ready),
    .io_deq_valid(cache_in_Q_io_deq_valid),
    .io_deq_bits_addr(cache_in_Q_io_deq_bits_addr),
    .io_deq_bits_inst(cache_in_Q_io_deq_bits_inst),
    .io_deq_bits_data(cache_in_Q_io_deq_bits_data),
    .io_deq_bits_src(cache_in_Q_io_deq_bits_src),
    .io_deq_bits_dst(cache_in_Q_io_deq_bits_dst),
    .io_deq_bits_msgType(cache_in_Q_io_deq_bits_msgType)
  );
  Queue_1 cache_out_Q ( // @[Router.scala 20:27]
    .clock(cache_out_Q_clock),
    .reset(cache_out_Q_reset),
    .io_enq_ready(cache_out_Q_io_enq_ready),
    .io_enq_valid(cache_out_Q_io_enq_valid),
    .io_enq_bits_addr(cache_out_Q_io_enq_bits_addr),
    .io_enq_bits_inst(cache_out_Q_io_enq_bits_inst),
    .io_enq_bits_data(cache_out_Q_io_enq_bits_data),
    .io_enq_bits_src(cache_out_Q_io_enq_bits_src),
    .io_enq_bits_dst(cache_out_Q_io_enq_bits_dst),
    .io_enq_bits_msgType(cache_out_Q_io_enq_bits_msgType),
    .io_deq_ready(cache_out_Q_io_deq_ready),
    .io_deq_valid(cache_out_Q_io_deq_valid),
    .io_deq_bits_addr(cache_out_Q_io_deq_bits_addr),
    .io_deq_bits_inst(cache_out_Q_io_deq_bits_inst),
    .io_deq_bits_data(cache_out_Q_io_deq_bits_data),
    .io_deq_bits_src(cache_out_Q_io_deq_bits_src),
    .io_deq_bits_dst(cache_out_Q_io_deq_bits_dst),
    .io_deq_bits_msgType(cache_out_Q_io_deq_bits_msgType)
  );
  Queue_3 in_Q ( // @[Router.scala 21:20]
    .clock(in_Q_clock),
    .reset(in_Q_reset),
    .io_enq_ready(in_Q_io_enq_ready),
    .io_enq_valid(in_Q_io_enq_valid),
    .io_enq_bits_addr(in_Q_io_enq_bits_addr),
    .io_enq_bits_inst(in_Q_io_enq_bits_inst),
    .io_enq_bits_data(in_Q_io_enq_bits_data),
    .io_enq_bits_src(in_Q_io_enq_bits_src),
    .io_enq_bits_dst(in_Q_io_enq_bits_dst),
    .io_enq_bits_msgType(in_Q_io_enq_bits_msgType),
    .io_deq_ready(in_Q_io_deq_ready),
    .io_deq_valid(in_Q_io_deq_valid),
    .io_deq_bits_addr(in_Q_io_deq_bits_addr),
    .io_deq_bits_inst(in_Q_io_deq_bits_inst),
    .io_deq_bits_data(in_Q_io_deq_bits_data),
    .io_deq_bits_src(in_Q_io_deq_bits_src),
    .io_deq_bits_dst(in_Q_io_deq_bits_dst),
    .io_deq_bits_msgType(in_Q_io_deq_bits_msgType)
  );
  RRArbiter arbiter ( // @[Router.scala 23:23]
    .clock(arbiter_clock),
    .io_in_0_ready(arbiter_io_in_0_ready),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_addr(arbiter_io_in_0_bits_addr),
    .io_in_0_bits_inst(arbiter_io_in_0_bits_inst),
    .io_in_0_bits_data(arbiter_io_in_0_bits_data),
    .io_in_0_bits_src(arbiter_io_in_0_bits_src),
    .io_in_0_bits_dst(arbiter_io_in_0_bits_dst),
    .io_in_0_bits_msgType(arbiter_io_in_0_bits_msgType),
    .io_in_1_ready(arbiter_io_in_1_ready),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_addr(arbiter_io_in_1_bits_addr),
    .io_in_1_bits_inst(arbiter_io_in_1_bits_inst),
    .io_in_1_bits_data(arbiter_io_in_1_bits_data),
    .io_in_1_bits_src(arbiter_io_in_1_bits_src),
    .io_in_1_bits_dst(arbiter_io_in_1_bits_dst),
    .io_in_1_bits_msgType(arbiter_io_in_1_bits_msgType),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_addr(arbiter_io_out_bits_addr),
    .io_out_bits_inst(arbiter_io_out_bits_inst),
    .io_out_bits_data(arbiter_io_out_bits_data),
    .io_out_bits_src(arbiter_io_out_bits_src),
    .io_out_bits_dst(arbiter_io_out_bits_dst),
    .io_out_bits_msgType(arbiter_io_out_bits_msgType),
    .io_chosen(arbiter_io_chosen)
  );
  assign io_cacheIn_ready = cache_in_Q_io_enq_ready; // @[Router.scala 25:21]
  assign io_cacheOut_valid = cache_out_Q_io_deq_valid; // @[Router.scala 26:15]
  assign io_cacheOut_bits_addr = cache_out_Q_io_deq_bits_addr; // @[Router.scala 26:15]
  assign io_cacheOut_bits_inst = cache_out_Q_io_deq_bits_inst; // @[Router.scala 26:15]
  assign io_cacheOut_bits_data = cache_out_Q_io_deq_bits_data; // @[Router.scala 26:15]
  assign io_cacheOut_bits_src = cache_out_Q_io_deq_bits_src; // @[Router.scala 26:15]
  assign io_in_ready = in_Q_io_enq_ready; // @[Router.scala 27:15]
  assign io_out_valid = arbiter_io_out_valid; // @[Router.scala 29:10]
  assign io_out_bits_addr = arbiter_io_out_bits_addr; // @[Router.scala 29:10]
  assign io_out_bits_inst = arbiter_io_out_bits_inst; // @[Router.scala 29:10]
  assign io_out_bits_data = arbiter_io_out_bits_data; // @[Router.scala 29:10]
  assign io_out_bits_src = arbiter_io_out_bits_src; // @[Router.scala 29:10]
  assign io_out_bits_dst = arbiter_io_out_bits_dst; // @[Router.scala 29:10]
  assign io_out_bits_msgType = arbiter_io_out_bits_msgType; // @[Router.scala 29:10]
  assign cache_in_Q_clock = clock;
  assign cache_in_Q_reset = reset;
  assign cache_in_Q_io_enq_valid = io_cacheIn_valid; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_addr = io_cacheIn_bits_addr; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_inst = 8'h2; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_data = io_cacheIn_bits_data; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_src = 3'h1; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_dst = io_cacheIn_bits_dst; // @[Router.scala 25:21]
  assign cache_in_Q_io_enq_bits_msgType = 2'h0; // @[Router.scala 25:21]
  assign cache_in_Q_io_deq_ready = arbiter_io_in_0_ready; // @[Router.scala 31:20]
  assign cache_out_Q_clock = clock;
  assign cache_out_Q_reset = reset;
  assign cache_out_Q_io_enq_valid = in_Q_io_deq_valid & _T; // @[Router.scala 34:28]
  assign cache_out_Q_io_enq_bits_addr = in_Q_io_deq_bits_addr; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_inst = in_Q_io_deq_bits_inst; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_data = in_Q_io_deq_bits_data; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_src = in_Q_io_deq_bits_src; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_dst = in_Q_io_deq_bits_dst; // @[Router.scala 33:27]
  assign cache_out_Q_io_enq_bits_msgType = in_Q_io_deq_bits_msgType; // @[Router.scala 33:27]
  assign cache_out_Q_io_deq_ready = io_cacheOut_ready; // @[Router.scala 26:15]
  assign in_Q_clock = clock;
  assign in_Q_reset = reset;
  assign in_Q_io_enq_valid = io_in_valid; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_addr = io_in_bits_addr; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_inst = io_in_bits_inst; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_data = io_in_bits_data; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_src = io_in_bits_src; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_dst = io_in_bits_dst; // @[Router.scala 27:15]
  assign in_Q_io_enq_bits_msgType = io_in_bits_msgType; // @[Router.scala 27:15]
  assign in_Q_io_deq_ready = _T_5 | _T_7; // @[Router.scala 38:21]
  assign arbiter_clock = clock;
  assign arbiter_io_in_0_valid = cache_in_Q_io_deq_valid; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_addr = cache_in_Q_io_deq_bits_addr; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_inst = cache_in_Q_io_deq_bits_inst; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_data = cache_in_Q_io_deq_bits_data; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_src = cache_in_Q_io_deq_bits_src; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_dst = cache_in_Q_io_deq_bits_dst; // @[Router.scala 31:20]
  assign arbiter_io_in_0_bits_msgType = cache_in_Q_io_deq_bits_msgType; // @[Router.scala 31:20]
  assign arbiter_io_in_1_valid = in_Q_io_deq_valid & _T_2; // @[Router.scala 37:26]
  assign arbiter_io_in_1_bits_addr = in_Q_io_deq_bits_addr; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_inst = in_Q_io_deq_bits_inst; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_data = in_Q_io_deq_bits_data; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_src = in_Q_io_deq_bits_src; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_dst = in_Q_io_deq_bits_dst; // @[Router.scala 36:25]
  assign arbiter_io_in_1_bits_msgType = in_Q_io_deq_bits_msgType; // @[Router.scala 36:25]
  assign arbiter_io_out_ready = io_out_ready; // @[Router.scala 29:10]
endmodule
module bipassLD(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [3:0]  io_in_bits_way,
  output        io_dataMem_in_valid,
  output [31:0] io_dataMem_in_bits_address,
  input  [63:0] io_dataMem_outputValue_0,
  output        io_out_valid,
  output [63:0] io_out_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [5:0] set = io_in_bits_addr[8:3]; // @[Gem5CacheLogic.scala 95:19]
  reg [63:0] dataRead_0; // @[elements.scala 323:27]
  wire [8:0] _T_1 = set * 6'h4; // @[elements.scala 327:39]
  wire [8:0] _GEN_0 = {{5'd0}, io_in_bits_way}; // @[elements.scala 327:49]
  wire [8:0] _T_3 = _T_1 + _GEN_0; // @[elements.scala 327:49]
  reg  _T_4; // @[elements.scala 331:28]
  assign io_dataMem_in_valid = io_in_valid; // @[elements.scala 325:25]
  assign io_dataMem_in_bits_address = {{23'd0}, _T_3}; // @[elements.scala 327:32]
  assign io_out_valid = _T_4; // @[elements.scala 331:18]
  assign io_out_bits_data = dataRead_0; // @[elements.scala 332:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  dataRead_0 = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  _T_4 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      dataRead_0 <= 64'h0;
    end else begin
      dataRead_0 <= io_dataMem_outputValue_0;
    end
    _T_4 <= io_in_valid;
  end
endmodule
module MemBank(
  input         clock,
  input         io_read_in_valid,
  input  [31:0] io_read_in_bits_address,
  output [63:0] io_read_outputValue_0,
  input         io_write_valid,
  input  [31:0] io_write_bits_address,
  input  [63:0] io_write_bits_inputValue_0
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [63:0] mems_0 [0:255]; // @[BankedMemory.scala 40:8]
  wire [63:0] mems_0__T_1_data; // @[BankedMemory.scala 40:8]
  wire [7:0] mems_0__T_1_addr; // @[BankedMemory.scala 40:8]
  wire [63:0] mems_0__T_5_data; // @[BankedMemory.scala 40:8]
  wire [7:0] mems_0__T_5_addr; // @[BankedMemory.scala 40:8]
  wire  mems_0__T_5_mask; // @[BankedMemory.scala 40:8]
  wire  mems_0__T_5_en; // @[BankedMemory.scala 40:8]
  assign mems_0__T_1_addr = io_read_in_bits_address[7:0];
  assign mems_0__T_1_data = mems_0[mems_0__T_1_addr]; // @[BankedMemory.scala 40:8]
  assign mems_0__T_5_data = io_write_bits_inputValue_0;
  assign mems_0__T_5_addr = io_write_bits_address[7:0];
  assign mems_0__T_5_mask = 1'h1;
  assign mems_0__T_5_en = io_write_valid;
  assign io_read_outputValue_0 = mems_0__T_1_data; // @[BankedMemory.scala 46:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mems_0[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mems_0__T_5_en & mems_0__T_5_mask) begin
      mems_0[mems_0__T_5_addr] <= mems_0__T_5_data; // @[BankedMemory.scala 40:8]
    end
  end
endmodule
module MemBank_1(
  input         clock,
  input         io_read_in_valid,
  input  [5:0]  io_read_in_bits_address,
  output [22:0] io_read_outputValue_0_tag,
  output [22:0] io_read_outputValue_1_tag,
  output [22:0] io_read_outputValue_2_tag,
  output [22:0] io_read_outputValue_3_tag,
  input         io_write_valid,
  input  [3:0]  io_write_bits_bank,
  input  [5:0]  io_write_bits_address,
  input  [22:0] io_write_bits_inputValue_0_tag,
  input  [22:0] io_write_bits_inputValue_1_tag,
  input  [22:0] io_write_bits_inputValue_2_tag,
  input  [22:0] io_write_bits_inputValue_3_tag
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
  reg [22:0] mems_0_tag [0:63]; // @[BankedMemory.scala 40:8]
  wire [22:0] mems_0_tag__T_data; // @[BankedMemory.scala 40:8]
  wire [5:0] mems_0_tag__T_addr; // @[BankedMemory.scala 40:8]
  wire [22:0] mems_0_tag__T_9_data; // @[BankedMemory.scala 40:8]
  wire [5:0] mems_0_tag__T_9_addr; // @[BankedMemory.scala 40:8]
  wire  mems_0_tag__T_9_mask; // @[BankedMemory.scala 40:8]
  wire  mems_0_tag__T_9_en; // @[BankedMemory.scala 40:8]
  reg [22:0] mems_1_tag [0:63]; // @[BankedMemory.scala 40:8]
  wire [22:0] mems_1_tag__T_1_data; // @[BankedMemory.scala 40:8]
  wire [5:0] mems_1_tag__T_1_addr; // @[BankedMemory.scala 40:8]
  wire [22:0] mems_1_tag__T_15_data; // @[BankedMemory.scala 40:8]
  wire [5:0] mems_1_tag__T_15_addr; // @[BankedMemory.scala 40:8]
  wire  mems_1_tag__T_15_mask; // @[BankedMemory.scala 40:8]
  wire  mems_1_tag__T_15_en; // @[BankedMemory.scala 40:8]
  reg [22:0] mems_2_tag [0:63]; // @[BankedMemory.scala 40:8]
  wire [22:0] mems_2_tag__T_2_data; // @[BankedMemory.scala 40:8]
  wire [5:0] mems_2_tag__T_2_addr; // @[BankedMemory.scala 40:8]
  wire [22:0] mems_2_tag__T_21_data; // @[BankedMemory.scala 40:8]
  wire [5:0] mems_2_tag__T_21_addr; // @[BankedMemory.scala 40:8]
  wire  mems_2_tag__T_21_mask; // @[BankedMemory.scala 40:8]
  wire  mems_2_tag__T_21_en; // @[BankedMemory.scala 40:8]
  reg [22:0] mems_3_tag [0:63]; // @[BankedMemory.scala 40:8]
  wire [22:0] mems_3_tag__T_3_data; // @[BankedMemory.scala 40:8]
  wire [5:0] mems_3_tag__T_3_addr; // @[BankedMemory.scala 40:8]
  wire [22:0] mems_3_tag__T_27_data; // @[BankedMemory.scala 40:8]
  wire [5:0] mems_3_tag__T_27_addr; // @[BankedMemory.scala 40:8]
  wire  mems_3_tag__T_27_mask; // @[BankedMemory.scala 40:8]
  wire  mems_3_tag__T_27_en; // @[BankedMemory.scala 40:8]
  wire  _GEN_19 = io_write_bits_bank[2] ? 1'h0 : io_write_bits_bank[3]; // @[BankedMemory.scala 57:82]
  wire  _GEN_29 = io_write_bits_bank[1] ? 1'h0 : io_write_bits_bank[2]; // @[BankedMemory.scala 57:82]
  wire  _GEN_34 = io_write_bits_bank[1] ? 1'h0 : _GEN_19; // @[BankedMemory.scala 57:82]
  wire  _GEN_44 = io_write_bits_bank[0] ? 1'h0 : io_write_bits_bank[1]; // @[BankedMemory.scala 57:82]
  wire  _GEN_49 = io_write_bits_bank[0] ? 1'h0 : _GEN_29; // @[BankedMemory.scala 57:82]
  wire  _GEN_54 = io_write_bits_bank[0] ? 1'h0 : _GEN_34; // @[BankedMemory.scala 57:82]
  assign mems_0_tag__T_addr = io_read_in_bits_address;
  assign mems_0_tag__T_data = mems_0_tag[mems_0_tag__T_addr]; // @[BankedMemory.scala 40:8]
  assign mems_0_tag__T_9_data = io_write_bits_inputValue_0_tag;
  assign mems_0_tag__T_9_addr = io_write_bits_address;
  assign mems_0_tag__T_9_mask = 1'h1;
  assign mems_0_tag__T_9_en = io_write_valid & io_write_bits_bank[0];
  assign mems_1_tag__T_1_addr = io_read_in_bits_address;
  assign mems_1_tag__T_1_data = mems_1_tag[mems_1_tag__T_1_addr]; // @[BankedMemory.scala 40:8]
  assign mems_1_tag__T_15_data = io_write_bits_inputValue_1_tag;
  assign mems_1_tag__T_15_addr = io_write_bits_address;
  assign mems_1_tag__T_15_mask = 1'h1;
  assign mems_1_tag__T_15_en = io_write_valid & _GEN_44;
  assign mems_2_tag__T_2_addr = io_read_in_bits_address;
  assign mems_2_tag__T_2_data = mems_2_tag[mems_2_tag__T_2_addr]; // @[BankedMemory.scala 40:8]
  assign mems_2_tag__T_21_data = io_write_bits_inputValue_2_tag;
  assign mems_2_tag__T_21_addr = io_write_bits_address;
  assign mems_2_tag__T_21_mask = 1'h1;
  assign mems_2_tag__T_21_en = io_write_valid & _GEN_49;
  assign mems_3_tag__T_3_addr = io_read_in_bits_address;
  assign mems_3_tag__T_3_data = mems_3_tag[mems_3_tag__T_3_addr]; // @[BankedMemory.scala 40:8]
  assign mems_3_tag__T_27_data = io_write_bits_inputValue_3_tag;
  assign mems_3_tag__T_27_addr = io_write_bits_address;
  assign mems_3_tag__T_27_mask = 1'h1;
  assign mems_3_tag__T_27_en = io_write_valid & _GEN_54;
  assign io_read_outputValue_0_tag = mems_0_tag__T_data; // @[BankedMemory.scala 46:42]
  assign io_read_outputValue_1_tag = mems_1_tag__T_1_data; // @[BankedMemory.scala 46:42]
  assign io_read_outputValue_2_tag = mems_2_tag__T_2_data; // @[BankedMemory.scala 46:42]
  assign io_read_outputValue_3_tag = mems_3_tag__T_3_data; // @[BankedMemory.scala 46:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    mems_0_tag[initvar] = _RAND_0[22:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    mems_1_tag[initvar] = _RAND_1[22:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    mems_2_tag[initvar] = _RAND_2[22:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    mems_3_tag[initvar] = _RAND_3[22:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mems_0_tag__T_9_en & mems_0_tag__T_9_mask) begin
      mems_0_tag[mems_0_tag__T_9_addr] <= mems_0_tag__T_9_data; // @[BankedMemory.scala 40:8]
    end
    if(mems_1_tag__T_15_en & mems_1_tag__T_15_mask) begin
      mems_1_tag[mems_1_tag__T_15_addr] <= mems_1_tag__T_15_data; // @[BankedMemory.scala 40:8]
    end
    if(mems_2_tag__T_21_en & mems_2_tag__T_21_mask) begin
      mems_2_tag[mems_2_tag__T_21_addr] <= mems_2_tag__T_21_data; // @[BankedMemory.scala 40:8]
    end
    if(mems_3_tag__T_27_en & mems_3_tag__T_27_mask) begin
      mems_3_tag[mems_3_tag__T_27_addr] <= mems_3_tag__T_27_data; // @[BankedMemory.scala 40:8]
    end
  end
endmodule
module Decoder(
  input  [27:0] io_inAction,
  output        io_outSignals_0,
  output        io_outSignals_1,
  output        io_outSignals_2,
  output        io_outSignals_3,
  output        io_outSignals_4,
  output        io_outSignals_5,
  output        io_outSignals_6,
  output        io_outSignals_7,
  output        io_outSignals_8
);
  assign io_outSignals_0 = io_inAction[0]; // @[elements.scala 21:19]
  assign io_outSignals_1 = io_inAction[1]; // @[elements.scala 21:19]
  assign io_outSignals_2 = io_inAction[2]; // @[elements.scala 21:19]
  assign io_outSignals_3 = io_inAction[3]; // @[elements.scala 21:19]
  assign io_outSignals_4 = io_inAction[4]; // @[elements.scala 21:19]
  assign io_outSignals_5 = io_inAction[5]; // @[elements.scala 21:19]
  assign io_outSignals_6 = io_inAction[6]; // @[elements.scala 21:19]
  assign io_outSignals_7 = io_inAction[7]; // @[elements.scala 21:19]
  assign io_outSignals_8 = io_inAction[8]; // @[elements.scala 21:19]
endmodule
module FindEmptyLine(
  input   io_data_0,
  input   io_data_1,
  input   io_data_2,
  input   io_data_3,
  output  io_value_valid
);
  wire  _T = ~io_data_0; // @[elements.scala 74:53]
  wire  _T_1 = ~io_data_1; // @[elements.scala 74:53]
  wire  _T_2 = ~io_data_2; // @[elements.scala 74:53]
  wire  _T_3 = ~io_data_3; // @[elements.scala 74:53]
  wire  _GEN_3 = _T_2 | _T_3; // @[elements.scala 74:66]
  wire  _GEN_5 = _T_1 | _GEN_3; // @[elements.scala 74:66]
  assign io_value_valid = _T | _GEN_5; // @[elements.scala 68:20 elements.scala 76:32 elements.scala 76:32 elements.scala 76:32 elements.scala 76:32]
endmodule
module Find(
  input  [22:0] io_key_tag,
  input  [22:0] io_data_0_tag,
  input  [22:0] io_data_1_tag,
  input  [22:0] io_data_2_tag,
  input  [22:0] io_data_3_tag,
  input         io_valid_0,
  input         io_valid_1,
  input         io_valid_2,
  input         io_valid_3,
  output        io_value_valid,
  output [31:0] io_value_bits
);
  wire  _T = io_data_0_tag == io_key_tag; // @[elements.scala 35:54]
  wire  _T_1 = io_data_1_tag == io_key_tag; // @[elements.scala 35:54]
  wire  _T_2 = io_data_2_tag == io_key_tag; // @[elements.scala 35:54]
  wire  _T_3 = io_data_3_tag == io_key_tag; // @[elements.scala 35:54]
  wire [3:0] bitmap = {_T_3,_T_2,_T_1,_T}; // @[Cat.scala 29:58]
  wire [3:0] _T_9 = {io_valid_3,io_valid_2,io_valid_1,io_valid_0}; // @[elements.scala 36:46]
  wire [3:0] _T_10 = bitmap & _T_9; // @[elements.scala 36:29]
  wire  _T_13 = |_T_10[3:2]; // @[OneHot.scala 32:14]
  wire [1:0] _T_14 = _T_10[3:2] | _T_10[1:0]; // @[OneHot.scala 32:28]
  wire [1:0] _T_16 = {_T_13,_T_14[1]}; // @[Cat.scala 29:58]
  assign io_value_valid = _T_10 != 4'h0; // @[elements.scala 39:20]
  assign io_value_bits = {{30'd0}, _T_16}; // @[elements.scala 38:19]
endmodule
module Gem5CacheLogic(
  input         clock,
  input         reset,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [63:0] io_cpu_req_bits_data,
  input  [27:0] io_cpu_req_bits_command,
  input  [2:0]  io_cpu_req_bits_way,
  input  [2:0]  io_cpu_req_bits_replaceWay,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_iswrite,
  output [2:0]  io_cpu_resp_bits_way,
  output        io_metaMem_write_valid,
  output [3:0]  io_metaMem_write_bits_bank,
  output [5:0]  io_metaMem_write_bits_address,
  output [22:0] io_metaMem_write_bits_inputValue_0_tag,
  output [22:0] io_metaMem_write_bits_inputValue_1_tag,
  output [22:0] io_metaMem_write_bits_inputValue_2_tag,
  output [22:0] io_metaMem_write_bits_inputValue_3_tag,
  output        io_dataMem_write_valid,
  output [31:0] io_dataMem_write_bits_address,
  output [63:0] io_dataMem_write_bits_inputValue_0,
  output        io_validTagBits_write_valid,
  output [63:0] io_validTagBits_write_bits_addr,
  output        io_validTagBits_write_bits_value,
  output        io_validTagBits_read_in_valid,
  output [63:0] io_validTagBits_read_in_bits_addr,
  input         io_validTagBits_read_out_0,
  input         io_validTagBits_read_out_1,
  input         io_validTagBits_read_out_2,
  input         io_validTagBits_read_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire [27:0] decoder_io_inAction; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_7; // @[Gem5CacheLogic.scala 188:23]
  wire  decoder_io_outSignals_8; // @[Gem5CacheLogic.scala 188:23]
  wire  emptyLine_io_data_0; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_data_1; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_data_2; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_data_3; // @[Gem5CacheLogic.scala 359:25]
  wire  emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 359:25]
  wire [22:0] tagFinder_io_key_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [22:0] tagFinder_io_data_0_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [22:0] tagFinder_io_data_1_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [22:0] tagFinder_io_data_2_tag; // @[Gem5CacheLogic.scala 362:25]
  wire [22:0] tagFinder_io_data_3_tag; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_0; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_1; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_2; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_valid_3; // @[Gem5CacheLogic.scala 362:25]
  wire  tagFinder_io_value_valid; // @[Gem5CacheLogic.scala 362:25]
  wire [31:0] tagFinder_io_value_bits; // @[Gem5CacheLogic.scala 362:25]
  reg [31:0] addr_reg; // @[Gem5CacheLogic.scala 202:25]
  reg [63:0] cpu_data; // @[Gem5CacheLogic.scala 203:25]
  reg [27:0] cpu_command; // @[Gem5CacheLogic.scala 205:28]
  reg [22:0] tag; // @[Gem5CacheLogic.scala 207:20]
  reg [5:0] set; // @[Gem5CacheLogic.scala 208:20]
  reg [3:0] wayInput; // @[Gem5CacheLogic.scala 209:25]
  reg [3:0] replaceWayInput; // @[Gem5CacheLogic.scala 210:32]
  wire  _T_3 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  wire [6:0] _GEN_53 = {{1'd0}, set}; // @[Gem5CacheLogic.scala 289:41]
  wire [12:0] _T_6 = _GEN_53 * 7'h40; // @[Gem5CacheLogic.scala 289:41]
  wire  signals_2 = decoder_io_outSignals_2; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  wayInvalid = wayInput == 4'h4; // @[Gem5CacheLogic.scala 351:27]
  wire  _T_28 = ~wayInvalid; // @[Gem5CacheLogic.scala 378:14]
  wire [3:0] _GEN_15 = _T_28 ? wayInput : 4'h4; // @[Gem5CacheLogic.scala 378:26]
  wire [3:0] way = signals_2 ? replaceWayInput : _GEN_15; // @[Gem5CacheLogic.scala 376:23]
  wire [12:0] _GEN_54 = {{9'd0}, way}; // @[Gem5CacheLogic.scala 289:51]
  wire [12:0] _T_8 = _T_6 + _GEN_54; // @[Gem5CacheLogic.scala 289:51]
  wire  signals_1 = decoder_io_outSignals_1; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_0 = decoder_io_outSignals_0; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_23 = signals_1 & signals_0; // @[Gem5CacheLogic.scala 367:37]
  wire  _T_24 = signals_2 | _T_23; // @[Gem5CacheLogic.scala 367:21]
  wire [8:0] _T_25 = set * 6'h4; // @[Gem5CacheLogic.scala 368:46]
  wire [8:0] _GEN_14 = _T_24 ? _T_25 : 9'h0; // @[Gem5CacheLogic.scala 367:53]
  wire [15:0] _T_29 = 16'h1 << way; // @[Gem5CacheLogic.scala 338:34]
  wire  signals_4 = decoder_io_outSignals_4; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_3 = decoder_io_outSignals_3; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire [8:0] _GEN_59 = {{5'd0}, way}; // @[Gem5CacheLogic.scala 403:50]
  wire [8:0] _T_44 = _T_25 + _GEN_59; // @[Gem5CacheLogic.scala 403:50]
  wire [31:0] _T_47 = tagFinder_io_value_valid ? tagFinder_io_value_bits : 32'h4; // @[Gem5CacheLogic.scala 424:25]
  wire [3:0] _GEN_45 = signals_2 ? way : 4'h4; // @[Gem5CacheLogic.scala 425:28]
  wire [31:0] _GEN_47 = _T_23 ? _T_47 : {{28'd0}, _GEN_45}; // @[Gem5CacheLogic.scala 423:39]
  wire  signals_5 = decoder_io_outSignals_5; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  signals_6 = decoder_io_outSignals_6; // @[Gem5CacheLogic.scala 228:21 Gem5CacheLogic.scala 299:11]
  wire  _T_52 = ~signals_6; // @[Gem5CacheLogic.scala 446:50]
  reg  _T_54; // @[Gem5CacheLogic.scala 455:38]
  reg  _T_57; // @[Gem5CacheLogic.scala 456:81]
  wire  _T_59 = ~emptyLine_io_value_valid; // @[Gem5CacheLogic.scala 460:26]
  wire  _T_60 = signals_2 & _T_59; // @[Gem5CacheLogic.scala 460:23]
  wire  _T_62 = ~reset; // @[Gem5CacheLogic.scala 461:13]
  wire [3:0] targetWayWire = _GEN_47[3:0]; // @[Gem5CacheLogic.scala 424:19 Gem5CacheLogic.scala 426:19]
  Decoder decoder ( // @[Gem5CacheLogic.scala 188:23]
    .io_inAction(decoder_io_inAction),
    .io_outSignals_0(decoder_io_outSignals_0),
    .io_outSignals_1(decoder_io_outSignals_1),
    .io_outSignals_2(decoder_io_outSignals_2),
    .io_outSignals_3(decoder_io_outSignals_3),
    .io_outSignals_4(decoder_io_outSignals_4),
    .io_outSignals_5(decoder_io_outSignals_5),
    .io_outSignals_6(decoder_io_outSignals_6),
    .io_outSignals_7(decoder_io_outSignals_7),
    .io_outSignals_8(decoder_io_outSignals_8)
  );
  FindEmptyLine emptyLine ( // @[Gem5CacheLogic.scala 359:25]
    .io_data_0(emptyLine_io_data_0),
    .io_data_1(emptyLine_io_data_1),
    .io_data_2(emptyLine_io_data_2),
    .io_data_3(emptyLine_io_data_3),
    .io_value_valid(emptyLine_io_value_valid)
  );
  Find tagFinder ( // @[Gem5CacheLogic.scala 362:25]
    .io_key_tag(tagFinder_io_key_tag),
    .io_data_0_tag(tagFinder_io_data_0_tag),
    .io_data_1_tag(tagFinder_io_data_1_tag),
    .io_data_2_tag(tagFinder_io_data_2_tag),
    .io_data_3_tag(tagFinder_io_data_3_tag),
    .io_valid_0(tagFinder_io_valid_0),
    .io_valid_1(tagFinder_io_valid_1),
    .io_valid_2(tagFinder_io_valid_2),
    .io_valid_3(tagFinder_io_valid_3),
    .io_value_valid(tagFinder_io_value_valid),
    .io_value_bits(tagFinder_io_value_bits)
  );
  assign io_cpu_req_ready = 1'h1; // @[Gem5CacheLogic.scala 302:20]
  assign io_cpu_resp_valid = _T_24 | _T_57; // @[Gem5CacheLogic.scala 456:24]
  assign io_cpu_resp_bits_iswrite = _T_54; // @[Gem5CacheLogic.scala 455:28]
  assign io_cpu_resp_bits_way = targetWayWire[2:0]; // @[Gem5CacheLogic.scala 453:24]
  assign io_metaMem_write_valid = signals_3 ? 1'h0 : signals_4; // @[Gem5CacheLogic.scala 346:26 Gem5CacheLogic.scala 330:19]
  assign io_metaMem_write_bits_bank = _T_29[3:0]; // @[Gem5CacheLogic.scala 338:27]
  assign io_metaMem_write_bits_address = set; // @[Gem5CacheLogic.scala 339:30]
  assign io_metaMem_write_bits_inputValue_0_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_metaMem_write_bits_inputValue_1_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_metaMem_write_bits_inputValue_2_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_metaMem_write_bits_inputValue_3_tag = tag; // @[Gem5CacheLogic.scala 418:45]
  assign io_dataMem_write_valid = decoder_io_outSignals_7; // @[Gem5CacheLogic.scala 347:26 Gem5CacheLogic.scala 330:19]
  assign io_dataMem_write_bits_address = {{19'd0}, _T_8}; // @[Gem5CacheLogic.scala 334:30]
  assign io_dataMem_write_bits_inputValue_0 = cpu_data; // @[Gem5CacheLogic.scala 397:38]
  assign io_validTagBits_write_valid = signals_5 | signals_6; // @[Gem5CacheLogic.scala 445:31]
  assign io_validTagBits_write_bits_addr = {{55'd0}, _T_44}; // @[Gem5CacheLogic.scala 444:35]
  assign io_validTagBits_write_bits_value = signals_5 | _T_52; // @[Gem5CacheLogic.scala 446:36]
  assign io_validTagBits_read_in_valid = signals_2 | _T_23; // @[Gem5CacheLogic.scala 373:33]
  assign io_validTagBits_read_in_bits_addr = {{55'd0}, _GEN_14}; // @[Gem5CacheLogic.scala 368:39 Gem5CacheLogic.scala 370:39]
  assign decoder_io_inAction = cpu_command; // @[Gem5CacheLogic.scala 298:23]
  assign emptyLine_io_data_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 360:21]
  assign emptyLine_io_data_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 360:21]
  assign emptyLine_io_data_2 = io_validTagBits_read_out_2; // @[Gem5CacheLogic.scala 360:21]
  assign emptyLine_io_data_3 = io_validTagBits_read_out_3; // @[Gem5CacheLogic.scala 360:21]
  assign tagFinder_io_key_tag = tag; // @[Gem5CacheLogic.scala 363:20]
  assign tagFinder_io_data_0_tag = 23'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_data_1_tag = 23'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_data_2_tag = 23'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_data_3_tag = 23'h0; // @[Gem5CacheLogic.scala 364:21]
  assign tagFinder_io_valid_0 = io_validTagBits_read_out_0; // @[Gem5CacheLogic.scala 365:22]
  assign tagFinder_io_valid_1 = io_validTagBits_read_out_1; // @[Gem5CacheLogic.scala 365:22]
  assign tagFinder_io_valid_2 = io_validTagBits_read_out_2; // @[Gem5CacheLogic.scala 365:22]
  assign tagFinder_io_valid_3 = io_validTagBits_read_out_3; // @[Gem5CacheLogic.scala 365:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  cpu_data = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  cpu_command = _RAND_2[27:0];
  _RAND_3 = {1{`RANDOM}};
  tag = _RAND_3[22:0];
  _RAND_4 = {1{`RANDOM}};
  set = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  wayInput = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  replaceWayInput = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  _T_54 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_57 = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr_reg <= 32'h0;
    end else if (_T_3) begin
      addr_reg <= io_cpu_req_bits_addr;
    end
    if (reset) begin
      cpu_data <= 64'h0;
    end else if (_T_3) begin
      cpu_data <= io_cpu_req_bits_data;
    end
    if (reset) begin
      cpu_command <= 28'h0;
    end else if (_T_3) begin
      cpu_command <= io_cpu_req_bits_command;
    end
    if (reset) begin
      tag <= 23'h0;
    end else if (_T_3) begin
      tag <= io_cpu_req_bits_addr[31:9];
    end
    if (reset) begin
      set <= 6'h0;
    end else if (_T_3) begin
      set <= io_cpu_req_bits_addr[8:3];
    end
    if (reset) begin
      wayInput <= 4'h4;
    end else if (_T_3) begin
      wayInput <= {{1'd0}, io_cpu_req_bits_way};
    end
    if (reset) begin
      replaceWayInput <= 4'h4;
    end else if (_T_3) begin
      replaceWayInput <= {{1'd0}, io_cpu_req_bits_replaceWay};
    end
    _T_54 <= decoder_io_outSignals_8;
    _T_57 <= decoder_io_outSignals_8;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_60 & _T_62) begin
          $fwrite(32'h80000002,"Replacement in Set: %d, Way: %d, Addr: %d\n",set,way,addr_reg); // @[Gem5CacheLogic.scala 461:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module FindMultiLine(
  input  [22:0] io_key_tag,
  input  [22:0] io_data_0_tag,
  input  [22:0] io_data_1_tag,
  input  [22:0] io_data_2_tag,
  input  [22:0] io_data_3_tag,
  output        io_value_bits_0,
  output        io_value_bits_1,
  output        io_value_bits_2,
  output        io_value_bits_3
);
  wire  _T = io_data_0_tag == io_key_tag; // @[elements.scala 54:54]
  wire  _T_1 = io_data_1_tag == io_key_tag; // @[elements.scala 54:54]
  wire  _T_2 = io_data_2_tag == io_key_tag; // @[elements.scala 54:54]
  wire  _T_3 = io_data_3_tag == io_key_tag; // @[elements.scala 54:54]
  wire [3:0] bitmap = {_T_3,_T_2,_T_1,_T}; // @[Cat.scala 29:58]
  assign io_value_bits_0 = bitmap[0]; // @[elements.scala 57:19]
  assign io_value_bits_1 = bitmap[1]; // @[elements.scala 57:19]
  assign io_value_bits_2 = bitmap[2]; // @[elements.scala 57:19]
  assign io_value_bits_3 = bitmap[3]; // @[elements.scala 57:19]
endmodule
module ProbeUnit(
  input         clock,
  input         reset,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [27:0] io_cpu_req_bits_command,
  output        io_cpu_resp_valid,
  output [2:0]  io_cpu_resp_bits_way,
  output        io_cpu_multiWay_valid,
  output [2:0]  io_cpu_multiWay_bits_way_0,
  output [2:0]  io_cpu_multiWay_bits_way_1,
  output [2:0]  io_cpu_multiWay_bits_way_2,
  output [2:0]  io_cpu_multiWay_bits_way_3,
  output [31:0] io_cpu_multiWay_bits_addr,
  output        io_metaMem_read_in_valid,
  output [5:0]  io_metaMem_read_in_bits_address,
  input  [22:0] io_metaMem_read_outputValue_0_tag,
  input  [22:0] io_metaMem_read_outputValue_1_tag,
  input  [22:0] io_metaMem_read_outputValue_2_tag,
  input  [22:0] io_metaMem_read_outputValue_3_tag,
  output        io_validTagBits_write_valid,
  output [63:0] io_validTagBits_write_bits_addr,
  output        io_validTagBits_write_bits_value,
  output        io_validTagBits_read_in_valid,
  output [63:0] io_validTagBits_read_in_bits_addr,
  input         io_validTagBits_read_out_0,
  input         io_validTagBits_read_out_1,
  input         io_validTagBits_read_out_2,
  input         io_validTagBits_read_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [27:0] decoder_io_inAction; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_0; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_1; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_2; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_3; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_4; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_5; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_6; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_7; // @[ProbeUnit.scala 48:23]
  wire  decoder_io_outSignals_8; // @[ProbeUnit.scala 48:23]
  wire  emptyLine_io_data_0; // @[ProbeUnit.scala 217:25]
  wire  emptyLine_io_data_1; // @[ProbeUnit.scala 217:25]
  wire  emptyLine_io_data_2; // @[ProbeUnit.scala 217:25]
  wire  emptyLine_io_data_3; // @[ProbeUnit.scala 217:25]
  wire  emptyLine_io_value_valid; // @[ProbeUnit.scala 217:25]
  wire [22:0] multiTagFinder_io_key_tag; // @[ProbeUnit.scala 220:30]
  wire [22:0] multiTagFinder_io_data_0_tag; // @[ProbeUnit.scala 220:30]
  wire [22:0] multiTagFinder_io_data_1_tag; // @[ProbeUnit.scala 220:30]
  wire [22:0] multiTagFinder_io_data_2_tag; // @[ProbeUnit.scala 220:30]
  wire [22:0] multiTagFinder_io_data_3_tag; // @[ProbeUnit.scala 220:30]
  wire  multiTagFinder_io_value_bits_0; // @[ProbeUnit.scala 220:30]
  wire  multiTagFinder_io_value_bits_1; // @[ProbeUnit.scala 220:30]
  wire  multiTagFinder_io_value_bits_2; // @[ProbeUnit.scala 220:30]
  wire  multiTagFinder_io_value_bits_3; // @[ProbeUnit.scala 220:30]
  wire [22:0] tagFinder_io_key_tag; // @[ProbeUnit.scala 221:25]
  wire [22:0] tagFinder_io_data_0_tag; // @[ProbeUnit.scala 221:25]
  wire [22:0] tagFinder_io_data_1_tag; // @[ProbeUnit.scala 221:25]
  wire [22:0] tagFinder_io_data_2_tag; // @[ProbeUnit.scala 221:25]
  wire [22:0] tagFinder_io_data_3_tag; // @[ProbeUnit.scala 221:25]
  wire  tagFinder_io_valid_0; // @[ProbeUnit.scala 221:25]
  wire  tagFinder_io_valid_1; // @[ProbeUnit.scala 221:25]
  wire  tagFinder_io_valid_2; // @[ProbeUnit.scala 221:25]
  wire  tagFinder_io_valid_3; // @[ProbeUnit.scala 221:25]
  wire  tagFinder_io_value_valid; // @[ProbeUnit.scala 221:25]
  wire [31:0] tagFinder_io_value_bits; // @[ProbeUnit.scala 221:25]
  reg [31:0] addr_reg; // @[ProbeUnit.scala 61:25]
  reg [27:0] cpu_command; // @[ProbeUnit.scala 64:28]
  reg [22:0] tag; // @[ProbeUnit.scala 66:20]
  reg [5:0] set; // @[ProbeUnit.scala 67:20]
  reg [3:0] wayInput; // @[ProbeUnit.scala 68:25]
  reg [3:0] replaceWayInput; // @[ProbeUnit.scala 69:32]
  wire  _T_4 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  wire  signals_2 = decoder_io_outSignals_2; // @[ProbeUnit.scala 87:21 ProbeUnit.scala 156:11]
  wire  wayInvalid = wayInput == 4'h4; // @[ProbeUnit.scala 209:27]
  wire  _T_30 = ~wayInvalid; // @[ProbeUnit.scala 245:14]
  wire [3:0] _GEN_15 = _T_30 ? wayInput : 4'h4; // @[ProbeUnit.scala 245:26]
  wire [3:0] way = signals_2 ? replaceWayInput : _GEN_15; // @[ProbeUnit.scala 243:23]
  wire  signals_1 = decoder_io_outSignals_1; // @[ProbeUnit.scala 87:21 ProbeUnit.scala 156:11]
  wire  signals_0 = decoder_io_outSignals_0; // @[ProbeUnit.scala 87:21 ProbeUnit.scala 156:11]
  wire  _T_25 = signals_1 & signals_0; // @[ProbeUnit.scala 234:37]
  wire  _T_26 = signals_2 | _T_25; // @[ProbeUnit.scala 234:21]
  wire [8:0] _T_27 = set * 6'h4; // @[ProbeUnit.scala 235:46]
  wire [8:0] _GEN_14 = _T_26 ? _T_27 : 9'h0; // @[ProbeUnit.scala 234:53]
  wire [8:0] _GEN_61 = {{5'd0}, way}; // @[ProbeUnit.scala 270:50]
  wire [8:0] _T_46 = _T_27 + _GEN_61; // @[ProbeUnit.scala 270:50]
  wire [31:0] _T_49 = tagFinder_io_value_valid ? tagFinder_io_value_bits : 32'h4; // @[ProbeUnit.scala 287:25]
  wire [3:0] _GEN_45 = signals_2 ? way : 4'h4; // @[ProbeUnit.scala 288:28]
  wire [31:0] _GEN_46 = _T_25 ? _T_49 : {{28'd0}, _GEN_45}; // @[ProbeUnit.scala 286:39]
  wire  _T_51 = multiTagFinder_io_value_bits_0; // @[ProbeUnit.scala 294:74]
  wire [2:0] _T_52 = _T_51 ? 3'h0 : 3'h4; // @[ProbeUnit.scala 294:35]
  wire  _T_53 = multiTagFinder_io_value_bits_1; // @[ProbeUnit.scala 294:74]
  wire [2:0] _T_54 = _T_53 ? 3'h1 : 3'h4; // @[ProbeUnit.scala 294:35]
  wire  _T_55 = multiTagFinder_io_value_bits_2; // @[ProbeUnit.scala 294:74]
  wire [2:0] _T_56 = _T_55 ? 3'h2 : 3'h4; // @[ProbeUnit.scala 294:35]
  wire  _T_57 = multiTagFinder_io_value_bits_3; // @[ProbeUnit.scala 294:74]
  wire [2:0] _T_58 = _T_57 ? 3'h3 : 3'h4; // @[ProbeUnit.scala 294:35]
  wire  signals_5 = decoder_io_outSignals_5; // @[ProbeUnit.scala 87:21 ProbeUnit.scala 156:11]
  wire  signals_6 = decoder_io_outSignals_6; // @[ProbeUnit.scala 87:21 ProbeUnit.scala 156:11]
  wire  _T_63 = ~signals_6; // @[ProbeUnit.scala 311:50]
  wire [3:0] targetWayWire = _GEN_46[3:0]; // @[ProbeUnit.scala 287:19 ProbeUnit.scala 289:19]
  Decoder decoder ( // @[ProbeUnit.scala 48:23]
    .io_inAction(decoder_io_inAction),
    .io_outSignals_0(decoder_io_outSignals_0),
    .io_outSignals_1(decoder_io_outSignals_1),
    .io_outSignals_2(decoder_io_outSignals_2),
    .io_outSignals_3(decoder_io_outSignals_3),
    .io_outSignals_4(decoder_io_outSignals_4),
    .io_outSignals_5(decoder_io_outSignals_5),
    .io_outSignals_6(decoder_io_outSignals_6),
    .io_outSignals_7(decoder_io_outSignals_7),
    .io_outSignals_8(decoder_io_outSignals_8)
  );
  FindEmptyLine emptyLine ( // @[ProbeUnit.scala 217:25]
    .io_data_0(emptyLine_io_data_0),
    .io_data_1(emptyLine_io_data_1),
    .io_data_2(emptyLine_io_data_2),
    .io_data_3(emptyLine_io_data_3),
    .io_value_valid(emptyLine_io_value_valid)
  );
  FindMultiLine multiTagFinder ( // @[ProbeUnit.scala 220:30]
    .io_key_tag(multiTagFinder_io_key_tag),
    .io_data_0_tag(multiTagFinder_io_data_0_tag),
    .io_data_1_tag(multiTagFinder_io_data_1_tag),
    .io_data_2_tag(multiTagFinder_io_data_2_tag),
    .io_data_3_tag(multiTagFinder_io_data_3_tag),
    .io_value_bits_0(multiTagFinder_io_value_bits_0),
    .io_value_bits_1(multiTagFinder_io_value_bits_1),
    .io_value_bits_2(multiTagFinder_io_value_bits_2),
    .io_value_bits_3(multiTagFinder_io_value_bits_3)
  );
  Find tagFinder ( // @[ProbeUnit.scala 221:25]
    .io_key_tag(tagFinder_io_key_tag),
    .io_data_0_tag(tagFinder_io_data_0_tag),
    .io_data_1_tag(tagFinder_io_data_1_tag),
    .io_data_2_tag(tagFinder_io_data_2_tag),
    .io_data_3_tag(tagFinder_io_data_3_tag),
    .io_valid_0(tagFinder_io_valid_0),
    .io_valid_1(tagFinder_io_valid_1),
    .io_valid_2(tagFinder_io_valid_2),
    .io_valid_3(tagFinder_io_valid_3),
    .io_value_valid(tagFinder_io_value_valid),
    .io_value_bits(tagFinder_io_value_bits)
  );
  assign io_cpu_req_ready = 1'h1; // @[ProbeUnit.scala 159:20]
  assign io_cpu_resp_valid = signals_1 & signals_0; // @[ProbeUnit.scala 321:24]
  assign io_cpu_resp_bits_way = targetWayWire[2:0]; // @[ProbeUnit.scala 318:24]
  assign io_cpu_multiWay_valid = io_cpu_resp_valid; // @[ProbeUnit.scala 322:25]
  assign io_cpu_multiWay_bits_way_0 = _T_25 ? _T_52 : 3'h0; // @[ProbeUnit.scala 315:28]
  assign io_cpu_multiWay_bits_way_1 = _T_25 ? _T_54 : 3'h0; // @[ProbeUnit.scala 315:28]
  assign io_cpu_multiWay_bits_way_2 = _T_25 ? _T_56 : 3'h0; // @[ProbeUnit.scala 315:28]
  assign io_cpu_multiWay_bits_way_3 = _T_25 ? _T_58 : 3'h0; // @[ProbeUnit.scala 315:28]
  assign io_cpu_multiWay_bits_addr = addr_reg; // @[ProbeUnit.scala 316:29]
  assign io_metaMem_read_in_valid = decoder_io_outSignals_3; // @[ProbeUnit.scala 206:28 ProbeUnit.scala 172:21]
  assign io_metaMem_read_in_bits_address = set; // @[ProbeUnit.scala 181:32]
  assign io_validTagBits_write_valid = signals_5 | signals_6; // @[ProbeUnit.scala 310:31]
  assign io_validTagBits_write_bits_addr = {{55'd0}, _T_46}; // @[ProbeUnit.scala 309:35]
  assign io_validTagBits_write_bits_value = signals_5 | _T_63; // @[ProbeUnit.scala 311:36]
  assign io_validTagBits_read_in_valid = signals_2 | _T_25; // @[ProbeUnit.scala 240:33]
  assign io_validTagBits_read_in_bits_addr = {{55'd0}, _GEN_14}; // @[ProbeUnit.scala 235:39 ProbeUnit.scala 237:39]
  assign decoder_io_inAction = cpu_command; // @[ProbeUnit.scala 155:23]
  assign emptyLine_io_data_0 = io_validTagBits_read_out_0; // @[ProbeUnit.scala 218:21]
  assign emptyLine_io_data_1 = io_validTagBits_read_out_1; // @[ProbeUnit.scala 218:21]
  assign emptyLine_io_data_2 = io_validTagBits_read_out_2; // @[ProbeUnit.scala 218:21]
  assign emptyLine_io_data_3 = io_validTagBits_read_out_3; // @[ProbeUnit.scala 218:21]
  assign multiTagFinder_io_key_tag = tag; // @[ProbeUnit.scala 227:25]
  assign multiTagFinder_io_data_0_tag = io_metaMem_read_outputValue_0_tag; // @[ProbeUnit.scala 228:26]
  assign multiTagFinder_io_data_1_tag = io_metaMem_read_outputValue_1_tag; // @[ProbeUnit.scala 228:26]
  assign multiTagFinder_io_data_2_tag = io_metaMem_read_outputValue_2_tag; // @[ProbeUnit.scala 228:26]
  assign multiTagFinder_io_data_3_tag = io_metaMem_read_outputValue_3_tag; // @[ProbeUnit.scala 228:26]
  assign tagFinder_io_key_tag = tag; // @[ProbeUnit.scala 223:20]
  assign tagFinder_io_data_0_tag = io_metaMem_read_outputValue_0_tag; // @[ProbeUnit.scala 224:21]
  assign tagFinder_io_data_1_tag = io_metaMem_read_outputValue_1_tag; // @[ProbeUnit.scala 224:21]
  assign tagFinder_io_data_2_tag = io_metaMem_read_outputValue_2_tag; // @[ProbeUnit.scala 224:21]
  assign tagFinder_io_data_3_tag = io_metaMem_read_outputValue_3_tag; // @[ProbeUnit.scala 224:21]
  assign tagFinder_io_valid_0 = io_validTagBits_read_out_0; // @[ProbeUnit.scala 225:22]
  assign tagFinder_io_valid_1 = io_validTagBits_read_out_1; // @[ProbeUnit.scala 225:22]
  assign tagFinder_io_valid_2 = io_validTagBits_read_out_2; // @[ProbeUnit.scala 225:22]
  assign tagFinder_io_valid_3 = io_validTagBits_read_out_3; // @[ProbeUnit.scala 225:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cpu_command = _RAND_1[27:0];
  _RAND_2 = {1{`RANDOM}};
  tag = _RAND_2[22:0];
  _RAND_3 = {1{`RANDOM}};
  set = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  wayInput = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  replaceWayInput = _RAND_5[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr_reg <= 32'h0;
    end else if (_T_4) begin
      addr_reg <= io_cpu_req_bits_addr;
    end
    if (reset) begin
      cpu_command <= 28'h0;
    end else if (_T_4) begin
      cpu_command <= io_cpu_req_bits_command;
    end else begin
      cpu_command <= 28'h0;
    end
    if (reset) begin
      tag <= 23'h0;
    end else if (_T_4) begin
      tag <= io_cpu_req_bits_addr[31:9];
    end
    if (reset) begin
      set <= 6'h0;
    end else if (_T_4) begin
      set <= io_cpu_req_bits_addr[8:3];
    end
    if (reset) begin
      wayInput <= 4'h4;
    end else if (_T_4) begin
      wayInput <= 4'h0;
    end
    if (reset) begin
      replaceWayInput <= 4'h4;
    end else if (_T_4) begin
      replaceWayInput <= 4'h0;
    end
  end
endmodule
module paralReg_1(
  input         clock,
  input         reset,
  input         io_port_0_write_valid,
  input  [63:0] io_port_0_write_bits_addr,
  input         io_port_0_write_bits_value,
  input         io_port_0_read_in_valid,
  input  [63:0] io_port_0_read_in_bits_addr,
  output        io_port_0_read_out_0,
  output        io_port_0_read_out_1,
  output        io_port_0_read_out_2,
  output        io_port_0_read_out_3,
  input         io_port_1_write_valid,
  input  [63:0] io_port_1_write_bits_addr,
  input         io_port_1_write_bits_value,
  input         io_port_1_read_in_valid,
  input  [63:0] io_port_1_read_in_bits_addr,
  output        io_port_1_read_out_0,
  output        io_port_1_read_out_1,
  output        io_port_1_read_out_2,
  output        io_port_1_read_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
`endif // RANDOMIZE_REG_INIT
  reg  content_0; // @[elements.scala 107:26]
  reg  content_1; // @[elements.scala 107:26]
  reg  content_2; // @[elements.scala 107:26]
  reg  content_3; // @[elements.scala 107:26]
  reg  content_4; // @[elements.scala 107:26]
  reg  content_5; // @[elements.scala 107:26]
  reg  content_6; // @[elements.scala 107:26]
  reg  content_7; // @[elements.scala 107:26]
  reg  content_8; // @[elements.scala 107:26]
  reg  content_9; // @[elements.scala 107:26]
  reg  content_10; // @[elements.scala 107:26]
  reg  content_11; // @[elements.scala 107:26]
  reg  content_12; // @[elements.scala 107:26]
  reg  content_13; // @[elements.scala 107:26]
  reg  content_14; // @[elements.scala 107:26]
  reg  content_15; // @[elements.scala 107:26]
  reg  content_16; // @[elements.scala 107:26]
  reg  content_17; // @[elements.scala 107:26]
  reg  content_18; // @[elements.scala 107:26]
  reg  content_19; // @[elements.scala 107:26]
  reg  content_20; // @[elements.scala 107:26]
  reg  content_21; // @[elements.scala 107:26]
  reg  content_22; // @[elements.scala 107:26]
  reg  content_23; // @[elements.scala 107:26]
  reg  content_24; // @[elements.scala 107:26]
  reg  content_25; // @[elements.scala 107:26]
  reg  content_26; // @[elements.scala 107:26]
  reg  content_27; // @[elements.scala 107:26]
  reg  content_28; // @[elements.scala 107:26]
  reg  content_29; // @[elements.scala 107:26]
  reg  content_30; // @[elements.scala 107:26]
  reg  content_31; // @[elements.scala 107:26]
  reg  content_32; // @[elements.scala 107:26]
  reg  content_33; // @[elements.scala 107:26]
  reg  content_34; // @[elements.scala 107:26]
  reg  content_35; // @[elements.scala 107:26]
  reg  content_36; // @[elements.scala 107:26]
  reg  content_37; // @[elements.scala 107:26]
  reg  content_38; // @[elements.scala 107:26]
  reg  content_39; // @[elements.scala 107:26]
  reg  content_40; // @[elements.scala 107:26]
  reg  content_41; // @[elements.scala 107:26]
  reg  content_42; // @[elements.scala 107:26]
  reg  content_43; // @[elements.scala 107:26]
  reg  content_44; // @[elements.scala 107:26]
  reg  content_45; // @[elements.scala 107:26]
  reg  content_46; // @[elements.scala 107:26]
  reg  content_47; // @[elements.scala 107:26]
  reg  content_48; // @[elements.scala 107:26]
  reg  content_49; // @[elements.scala 107:26]
  reg  content_50; // @[elements.scala 107:26]
  reg  content_51; // @[elements.scala 107:26]
  reg  content_52; // @[elements.scala 107:26]
  reg  content_53; // @[elements.scala 107:26]
  reg  content_54; // @[elements.scala 107:26]
  reg  content_55; // @[elements.scala 107:26]
  reg  content_56; // @[elements.scala 107:26]
  reg  content_57; // @[elements.scala 107:26]
  reg  content_58; // @[elements.scala 107:26]
  reg  content_59; // @[elements.scala 107:26]
  reg  content_60; // @[elements.scala 107:26]
  reg  content_61; // @[elements.scala 107:26]
  reg  content_62; // @[elements.scala 107:26]
  reg  content_63; // @[elements.scala 107:26]
  reg  content_64; // @[elements.scala 107:26]
  reg  content_65; // @[elements.scala 107:26]
  reg  content_66; // @[elements.scala 107:26]
  reg  content_67; // @[elements.scala 107:26]
  reg  content_68; // @[elements.scala 107:26]
  reg  content_69; // @[elements.scala 107:26]
  reg  content_70; // @[elements.scala 107:26]
  reg  content_71; // @[elements.scala 107:26]
  reg  content_72; // @[elements.scala 107:26]
  reg  content_73; // @[elements.scala 107:26]
  reg  content_74; // @[elements.scala 107:26]
  reg  content_75; // @[elements.scala 107:26]
  reg  content_76; // @[elements.scala 107:26]
  reg  content_77; // @[elements.scala 107:26]
  reg  content_78; // @[elements.scala 107:26]
  reg  content_79; // @[elements.scala 107:26]
  reg  content_80; // @[elements.scala 107:26]
  reg  content_81; // @[elements.scala 107:26]
  reg  content_82; // @[elements.scala 107:26]
  reg  content_83; // @[elements.scala 107:26]
  reg  content_84; // @[elements.scala 107:26]
  reg  content_85; // @[elements.scala 107:26]
  reg  content_86; // @[elements.scala 107:26]
  reg  content_87; // @[elements.scala 107:26]
  reg  content_88; // @[elements.scala 107:26]
  reg  content_89; // @[elements.scala 107:26]
  reg  content_90; // @[elements.scala 107:26]
  reg  content_91; // @[elements.scala 107:26]
  reg  content_92; // @[elements.scala 107:26]
  reg  content_93; // @[elements.scala 107:26]
  reg  content_94; // @[elements.scala 107:26]
  reg  content_95; // @[elements.scala 107:26]
  reg  content_96; // @[elements.scala 107:26]
  reg  content_97; // @[elements.scala 107:26]
  reg  content_98; // @[elements.scala 107:26]
  reg  content_99; // @[elements.scala 107:26]
  reg  content_100; // @[elements.scala 107:26]
  reg  content_101; // @[elements.scala 107:26]
  reg  content_102; // @[elements.scala 107:26]
  reg  content_103; // @[elements.scala 107:26]
  reg  content_104; // @[elements.scala 107:26]
  reg  content_105; // @[elements.scala 107:26]
  reg  content_106; // @[elements.scala 107:26]
  reg  content_107; // @[elements.scala 107:26]
  reg  content_108; // @[elements.scala 107:26]
  reg  content_109; // @[elements.scala 107:26]
  reg  content_110; // @[elements.scala 107:26]
  reg  content_111; // @[elements.scala 107:26]
  reg  content_112; // @[elements.scala 107:26]
  reg  content_113; // @[elements.scala 107:26]
  reg  content_114; // @[elements.scala 107:26]
  reg  content_115; // @[elements.scala 107:26]
  reg  content_116; // @[elements.scala 107:26]
  reg  content_117; // @[elements.scala 107:26]
  reg  content_118; // @[elements.scala 107:26]
  reg  content_119; // @[elements.scala 107:26]
  reg  content_120; // @[elements.scala 107:26]
  reg  content_121; // @[elements.scala 107:26]
  reg  content_122; // @[elements.scala 107:26]
  reg  content_123; // @[elements.scala 107:26]
  reg  content_124; // @[elements.scala 107:26]
  reg  content_125; // @[elements.scala 107:26]
  reg  content_126; // @[elements.scala 107:26]
  reg  content_127; // @[elements.scala 107:26]
  reg  content_128; // @[elements.scala 107:26]
  reg  content_129; // @[elements.scala 107:26]
  reg  content_130; // @[elements.scala 107:26]
  reg  content_131; // @[elements.scala 107:26]
  reg  content_132; // @[elements.scala 107:26]
  reg  content_133; // @[elements.scala 107:26]
  reg  content_134; // @[elements.scala 107:26]
  reg  content_135; // @[elements.scala 107:26]
  reg  content_136; // @[elements.scala 107:26]
  reg  content_137; // @[elements.scala 107:26]
  reg  content_138; // @[elements.scala 107:26]
  reg  content_139; // @[elements.scala 107:26]
  reg  content_140; // @[elements.scala 107:26]
  reg  content_141; // @[elements.scala 107:26]
  reg  content_142; // @[elements.scala 107:26]
  reg  content_143; // @[elements.scala 107:26]
  reg  content_144; // @[elements.scala 107:26]
  reg  content_145; // @[elements.scala 107:26]
  reg  content_146; // @[elements.scala 107:26]
  reg  content_147; // @[elements.scala 107:26]
  reg  content_148; // @[elements.scala 107:26]
  reg  content_149; // @[elements.scala 107:26]
  reg  content_150; // @[elements.scala 107:26]
  reg  content_151; // @[elements.scala 107:26]
  reg  content_152; // @[elements.scala 107:26]
  reg  content_153; // @[elements.scala 107:26]
  reg  content_154; // @[elements.scala 107:26]
  reg  content_155; // @[elements.scala 107:26]
  reg  content_156; // @[elements.scala 107:26]
  reg  content_157; // @[elements.scala 107:26]
  reg  content_158; // @[elements.scala 107:26]
  reg  content_159; // @[elements.scala 107:26]
  reg  content_160; // @[elements.scala 107:26]
  reg  content_161; // @[elements.scala 107:26]
  reg  content_162; // @[elements.scala 107:26]
  reg  content_163; // @[elements.scala 107:26]
  reg  content_164; // @[elements.scala 107:26]
  reg  content_165; // @[elements.scala 107:26]
  reg  content_166; // @[elements.scala 107:26]
  reg  content_167; // @[elements.scala 107:26]
  reg  content_168; // @[elements.scala 107:26]
  reg  content_169; // @[elements.scala 107:26]
  reg  content_170; // @[elements.scala 107:26]
  reg  content_171; // @[elements.scala 107:26]
  reg  content_172; // @[elements.scala 107:26]
  reg  content_173; // @[elements.scala 107:26]
  reg  content_174; // @[elements.scala 107:26]
  reg  content_175; // @[elements.scala 107:26]
  reg  content_176; // @[elements.scala 107:26]
  reg  content_177; // @[elements.scala 107:26]
  reg  content_178; // @[elements.scala 107:26]
  reg  content_179; // @[elements.scala 107:26]
  reg  content_180; // @[elements.scala 107:26]
  reg  content_181; // @[elements.scala 107:26]
  reg  content_182; // @[elements.scala 107:26]
  reg  content_183; // @[elements.scala 107:26]
  reg  content_184; // @[elements.scala 107:26]
  reg  content_185; // @[elements.scala 107:26]
  reg  content_186; // @[elements.scala 107:26]
  reg  content_187; // @[elements.scala 107:26]
  reg  content_188; // @[elements.scala 107:26]
  reg  content_189; // @[elements.scala 107:26]
  reg  content_190; // @[elements.scala 107:26]
  reg  content_191; // @[elements.scala 107:26]
  reg  content_192; // @[elements.scala 107:26]
  reg  content_193; // @[elements.scala 107:26]
  reg  content_194; // @[elements.scala 107:26]
  reg  content_195; // @[elements.scala 107:26]
  reg  content_196; // @[elements.scala 107:26]
  reg  content_197; // @[elements.scala 107:26]
  reg  content_198; // @[elements.scala 107:26]
  reg  content_199; // @[elements.scala 107:26]
  reg  content_200; // @[elements.scala 107:26]
  reg  content_201; // @[elements.scala 107:26]
  reg  content_202; // @[elements.scala 107:26]
  reg  content_203; // @[elements.scala 107:26]
  reg  content_204; // @[elements.scala 107:26]
  reg  content_205; // @[elements.scala 107:26]
  reg  content_206; // @[elements.scala 107:26]
  reg  content_207; // @[elements.scala 107:26]
  reg  content_208; // @[elements.scala 107:26]
  reg  content_209; // @[elements.scala 107:26]
  reg  content_210; // @[elements.scala 107:26]
  reg  content_211; // @[elements.scala 107:26]
  reg  content_212; // @[elements.scala 107:26]
  reg  content_213; // @[elements.scala 107:26]
  reg  content_214; // @[elements.scala 107:26]
  reg  content_215; // @[elements.scala 107:26]
  reg  content_216; // @[elements.scala 107:26]
  reg  content_217; // @[elements.scala 107:26]
  reg  content_218; // @[elements.scala 107:26]
  reg  content_219; // @[elements.scala 107:26]
  reg  content_220; // @[elements.scala 107:26]
  reg  content_221; // @[elements.scala 107:26]
  reg  content_222; // @[elements.scala 107:26]
  reg  content_223; // @[elements.scala 107:26]
  reg  content_224; // @[elements.scala 107:26]
  reg  content_225; // @[elements.scala 107:26]
  reg  content_226; // @[elements.scala 107:26]
  reg  content_227; // @[elements.scala 107:26]
  reg  content_228; // @[elements.scala 107:26]
  reg  content_229; // @[elements.scala 107:26]
  reg  content_230; // @[elements.scala 107:26]
  reg  content_231; // @[elements.scala 107:26]
  reg  content_232; // @[elements.scala 107:26]
  reg  content_233; // @[elements.scala 107:26]
  reg  content_234; // @[elements.scala 107:26]
  reg  content_235; // @[elements.scala 107:26]
  reg  content_236; // @[elements.scala 107:26]
  reg  content_237; // @[elements.scala 107:26]
  reg  content_238; // @[elements.scala 107:26]
  reg  content_239; // @[elements.scala 107:26]
  reg  content_240; // @[elements.scala 107:26]
  reg  content_241; // @[elements.scala 107:26]
  reg  content_242; // @[elements.scala 107:26]
  reg  content_243; // @[elements.scala 107:26]
  reg  content_244; // @[elements.scala 107:26]
  reg  content_245; // @[elements.scala 107:26]
  reg  content_246; // @[elements.scala 107:26]
  reg  content_247; // @[elements.scala 107:26]
  reg  content_248; // @[elements.scala 107:26]
  reg  content_249; // @[elements.scala 107:26]
  reg  content_250; // @[elements.scala 107:26]
  reg  content_251; // @[elements.scala 107:26]
  reg  content_252; // @[elements.scala 107:26]
  reg  content_253; // @[elements.scala 107:26]
  reg  content_254; // @[elements.scala 107:26]
  reg  content_255; // @[elements.scala 107:26]
  wire [64:0] _T_1 = {{1'd0}, io_port_0_read_in_bits_addr}; // @[elements.scala 118:104]
  wire [63:0] _T_5 = io_port_0_read_in_bits_addr + 64'h1; // @[elements.scala 118:104]
  wire [63:0] _T_8 = io_port_0_read_in_bits_addr + 64'h2; // @[elements.scala 118:104]
  wire [63:0] _T_11 = io_port_0_read_in_bits_addr + 64'h3; // @[elements.scala 118:104]
  wire  _GEN_1 = 8'h1 == _T_5[7:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_2 = 8'h2 == _T_5[7:0] ? content_2 : _GEN_1; // @[Cat.scala 29:58]
  wire  _GEN_3 = 8'h3 == _T_5[7:0] ? content_3 : _GEN_2; // @[Cat.scala 29:58]
  wire  _GEN_4 = 8'h4 == _T_5[7:0] ? content_4 : _GEN_3; // @[Cat.scala 29:58]
  wire  _GEN_5 = 8'h5 == _T_5[7:0] ? content_5 : _GEN_4; // @[Cat.scala 29:58]
  wire  _GEN_6 = 8'h6 == _T_5[7:0] ? content_6 : _GEN_5; // @[Cat.scala 29:58]
  wire  _GEN_7 = 8'h7 == _T_5[7:0] ? content_7 : _GEN_6; // @[Cat.scala 29:58]
  wire  _GEN_8 = 8'h8 == _T_5[7:0] ? content_8 : _GEN_7; // @[Cat.scala 29:58]
  wire  _GEN_9 = 8'h9 == _T_5[7:0] ? content_9 : _GEN_8; // @[Cat.scala 29:58]
  wire  _GEN_10 = 8'ha == _T_5[7:0] ? content_10 : _GEN_9; // @[Cat.scala 29:58]
  wire  _GEN_11 = 8'hb == _T_5[7:0] ? content_11 : _GEN_10; // @[Cat.scala 29:58]
  wire  _GEN_12 = 8'hc == _T_5[7:0] ? content_12 : _GEN_11; // @[Cat.scala 29:58]
  wire  _GEN_13 = 8'hd == _T_5[7:0] ? content_13 : _GEN_12; // @[Cat.scala 29:58]
  wire  _GEN_14 = 8'he == _T_5[7:0] ? content_14 : _GEN_13; // @[Cat.scala 29:58]
  wire  _GEN_15 = 8'hf == _T_5[7:0] ? content_15 : _GEN_14; // @[Cat.scala 29:58]
  wire  _GEN_16 = 8'h10 == _T_5[7:0] ? content_16 : _GEN_15; // @[Cat.scala 29:58]
  wire  _GEN_17 = 8'h11 == _T_5[7:0] ? content_17 : _GEN_16; // @[Cat.scala 29:58]
  wire  _GEN_18 = 8'h12 == _T_5[7:0] ? content_18 : _GEN_17; // @[Cat.scala 29:58]
  wire  _GEN_19 = 8'h13 == _T_5[7:0] ? content_19 : _GEN_18; // @[Cat.scala 29:58]
  wire  _GEN_20 = 8'h14 == _T_5[7:0] ? content_20 : _GEN_19; // @[Cat.scala 29:58]
  wire  _GEN_21 = 8'h15 == _T_5[7:0] ? content_21 : _GEN_20; // @[Cat.scala 29:58]
  wire  _GEN_22 = 8'h16 == _T_5[7:0] ? content_22 : _GEN_21; // @[Cat.scala 29:58]
  wire  _GEN_23 = 8'h17 == _T_5[7:0] ? content_23 : _GEN_22; // @[Cat.scala 29:58]
  wire  _GEN_24 = 8'h18 == _T_5[7:0] ? content_24 : _GEN_23; // @[Cat.scala 29:58]
  wire  _GEN_25 = 8'h19 == _T_5[7:0] ? content_25 : _GEN_24; // @[Cat.scala 29:58]
  wire  _GEN_26 = 8'h1a == _T_5[7:0] ? content_26 : _GEN_25; // @[Cat.scala 29:58]
  wire  _GEN_27 = 8'h1b == _T_5[7:0] ? content_27 : _GEN_26; // @[Cat.scala 29:58]
  wire  _GEN_28 = 8'h1c == _T_5[7:0] ? content_28 : _GEN_27; // @[Cat.scala 29:58]
  wire  _GEN_29 = 8'h1d == _T_5[7:0] ? content_29 : _GEN_28; // @[Cat.scala 29:58]
  wire  _GEN_30 = 8'h1e == _T_5[7:0] ? content_30 : _GEN_29; // @[Cat.scala 29:58]
  wire  _GEN_31 = 8'h1f == _T_5[7:0] ? content_31 : _GEN_30; // @[Cat.scala 29:58]
  wire  _GEN_32 = 8'h20 == _T_5[7:0] ? content_32 : _GEN_31; // @[Cat.scala 29:58]
  wire  _GEN_33 = 8'h21 == _T_5[7:0] ? content_33 : _GEN_32; // @[Cat.scala 29:58]
  wire  _GEN_34 = 8'h22 == _T_5[7:0] ? content_34 : _GEN_33; // @[Cat.scala 29:58]
  wire  _GEN_35 = 8'h23 == _T_5[7:0] ? content_35 : _GEN_34; // @[Cat.scala 29:58]
  wire  _GEN_36 = 8'h24 == _T_5[7:0] ? content_36 : _GEN_35; // @[Cat.scala 29:58]
  wire  _GEN_37 = 8'h25 == _T_5[7:0] ? content_37 : _GEN_36; // @[Cat.scala 29:58]
  wire  _GEN_38 = 8'h26 == _T_5[7:0] ? content_38 : _GEN_37; // @[Cat.scala 29:58]
  wire  _GEN_39 = 8'h27 == _T_5[7:0] ? content_39 : _GEN_38; // @[Cat.scala 29:58]
  wire  _GEN_40 = 8'h28 == _T_5[7:0] ? content_40 : _GEN_39; // @[Cat.scala 29:58]
  wire  _GEN_41 = 8'h29 == _T_5[7:0] ? content_41 : _GEN_40; // @[Cat.scala 29:58]
  wire  _GEN_42 = 8'h2a == _T_5[7:0] ? content_42 : _GEN_41; // @[Cat.scala 29:58]
  wire  _GEN_43 = 8'h2b == _T_5[7:0] ? content_43 : _GEN_42; // @[Cat.scala 29:58]
  wire  _GEN_44 = 8'h2c == _T_5[7:0] ? content_44 : _GEN_43; // @[Cat.scala 29:58]
  wire  _GEN_45 = 8'h2d == _T_5[7:0] ? content_45 : _GEN_44; // @[Cat.scala 29:58]
  wire  _GEN_46 = 8'h2e == _T_5[7:0] ? content_46 : _GEN_45; // @[Cat.scala 29:58]
  wire  _GEN_47 = 8'h2f == _T_5[7:0] ? content_47 : _GEN_46; // @[Cat.scala 29:58]
  wire  _GEN_48 = 8'h30 == _T_5[7:0] ? content_48 : _GEN_47; // @[Cat.scala 29:58]
  wire  _GEN_49 = 8'h31 == _T_5[7:0] ? content_49 : _GEN_48; // @[Cat.scala 29:58]
  wire  _GEN_50 = 8'h32 == _T_5[7:0] ? content_50 : _GEN_49; // @[Cat.scala 29:58]
  wire  _GEN_51 = 8'h33 == _T_5[7:0] ? content_51 : _GEN_50; // @[Cat.scala 29:58]
  wire  _GEN_52 = 8'h34 == _T_5[7:0] ? content_52 : _GEN_51; // @[Cat.scala 29:58]
  wire  _GEN_53 = 8'h35 == _T_5[7:0] ? content_53 : _GEN_52; // @[Cat.scala 29:58]
  wire  _GEN_54 = 8'h36 == _T_5[7:0] ? content_54 : _GEN_53; // @[Cat.scala 29:58]
  wire  _GEN_55 = 8'h37 == _T_5[7:0] ? content_55 : _GEN_54; // @[Cat.scala 29:58]
  wire  _GEN_56 = 8'h38 == _T_5[7:0] ? content_56 : _GEN_55; // @[Cat.scala 29:58]
  wire  _GEN_57 = 8'h39 == _T_5[7:0] ? content_57 : _GEN_56; // @[Cat.scala 29:58]
  wire  _GEN_58 = 8'h3a == _T_5[7:0] ? content_58 : _GEN_57; // @[Cat.scala 29:58]
  wire  _GEN_59 = 8'h3b == _T_5[7:0] ? content_59 : _GEN_58; // @[Cat.scala 29:58]
  wire  _GEN_60 = 8'h3c == _T_5[7:0] ? content_60 : _GEN_59; // @[Cat.scala 29:58]
  wire  _GEN_61 = 8'h3d == _T_5[7:0] ? content_61 : _GEN_60; // @[Cat.scala 29:58]
  wire  _GEN_62 = 8'h3e == _T_5[7:0] ? content_62 : _GEN_61; // @[Cat.scala 29:58]
  wire  _GEN_63 = 8'h3f == _T_5[7:0] ? content_63 : _GEN_62; // @[Cat.scala 29:58]
  wire  _GEN_64 = 8'h40 == _T_5[7:0] ? content_64 : _GEN_63; // @[Cat.scala 29:58]
  wire  _GEN_65 = 8'h41 == _T_5[7:0] ? content_65 : _GEN_64; // @[Cat.scala 29:58]
  wire  _GEN_66 = 8'h42 == _T_5[7:0] ? content_66 : _GEN_65; // @[Cat.scala 29:58]
  wire  _GEN_67 = 8'h43 == _T_5[7:0] ? content_67 : _GEN_66; // @[Cat.scala 29:58]
  wire  _GEN_68 = 8'h44 == _T_5[7:0] ? content_68 : _GEN_67; // @[Cat.scala 29:58]
  wire  _GEN_69 = 8'h45 == _T_5[7:0] ? content_69 : _GEN_68; // @[Cat.scala 29:58]
  wire  _GEN_70 = 8'h46 == _T_5[7:0] ? content_70 : _GEN_69; // @[Cat.scala 29:58]
  wire  _GEN_71 = 8'h47 == _T_5[7:0] ? content_71 : _GEN_70; // @[Cat.scala 29:58]
  wire  _GEN_72 = 8'h48 == _T_5[7:0] ? content_72 : _GEN_71; // @[Cat.scala 29:58]
  wire  _GEN_73 = 8'h49 == _T_5[7:0] ? content_73 : _GEN_72; // @[Cat.scala 29:58]
  wire  _GEN_74 = 8'h4a == _T_5[7:0] ? content_74 : _GEN_73; // @[Cat.scala 29:58]
  wire  _GEN_75 = 8'h4b == _T_5[7:0] ? content_75 : _GEN_74; // @[Cat.scala 29:58]
  wire  _GEN_76 = 8'h4c == _T_5[7:0] ? content_76 : _GEN_75; // @[Cat.scala 29:58]
  wire  _GEN_77 = 8'h4d == _T_5[7:0] ? content_77 : _GEN_76; // @[Cat.scala 29:58]
  wire  _GEN_78 = 8'h4e == _T_5[7:0] ? content_78 : _GEN_77; // @[Cat.scala 29:58]
  wire  _GEN_79 = 8'h4f == _T_5[7:0] ? content_79 : _GEN_78; // @[Cat.scala 29:58]
  wire  _GEN_80 = 8'h50 == _T_5[7:0] ? content_80 : _GEN_79; // @[Cat.scala 29:58]
  wire  _GEN_81 = 8'h51 == _T_5[7:0] ? content_81 : _GEN_80; // @[Cat.scala 29:58]
  wire  _GEN_82 = 8'h52 == _T_5[7:0] ? content_82 : _GEN_81; // @[Cat.scala 29:58]
  wire  _GEN_83 = 8'h53 == _T_5[7:0] ? content_83 : _GEN_82; // @[Cat.scala 29:58]
  wire  _GEN_84 = 8'h54 == _T_5[7:0] ? content_84 : _GEN_83; // @[Cat.scala 29:58]
  wire  _GEN_85 = 8'h55 == _T_5[7:0] ? content_85 : _GEN_84; // @[Cat.scala 29:58]
  wire  _GEN_86 = 8'h56 == _T_5[7:0] ? content_86 : _GEN_85; // @[Cat.scala 29:58]
  wire  _GEN_87 = 8'h57 == _T_5[7:0] ? content_87 : _GEN_86; // @[Cat.scala 29:58]
  wire  _GEN_88 = 8'h58 == _T_5[7:0] ? content_88 : _GEN_87; // @[Cat.scala 29:58]
  wire  _GEN_89 = 8'h59 == _T_5[7:0] ? content_89 : _GEN_88; // @[Cat.scala 29:58]
  wire  _GEN_90 = 8'h5a == _T_5[7:0] ? content_90 : _GEN_89; // @[Cat.scala 29:58]
  wire  _GEN_91 = 8'h5b == _T_5[7:0] ? content_91 : _GEN_90; // @[Cat.scala 29:58]
  wire  _GEN_92 = 8'h5c == _T_5[7:0] ? content_92 : _GEN_91; // @[Cat.scala 29:58]
  wire  _GEN_93 = 8'h5d == _T_5[7:0] ? content_93 : _GEN_92; // @[Cat.scala 29:58]
  wire  _GEN_94 = 8'h5e == _T_5[7:0] ? content_94 : _GEN_93; // @[Cat.scala 29:58]
  wire  _GEN_95 = 8'h5f == _T_5[7:0] ? content_95 : _GEN_94; // @[Cat.scala 29:58]
  wire  _GEN_96 = 8'h60 == _T_5[7:0] ? content_96 : _GEN_95; // @[Cat.scala 29:58]
  wire  _GEN_97 = 8'h61 == _T_5[7:0] ? content_97 : _GEN_96; // @[Cat.scala 29:58]
  wire  _GEN_98 = 8'h62 == _T_5[7:0] ? content_98 : _GEN_97; // @[Cat.scala 29:58]
  wire  _GEN_99 = 8'h63 == _T_5[7:0] ? content_99 : _GEN_98; // @[Cat.scala 29:58]
  wire  _GEN_100 = 8'h64 == _T_5[7:0] ? content_100 : _GEN_99; // @[Cat.scala 29:58]
  wire  _GEN_101 = 8'h65 == _T_5[7:0] ? content_101 : _GEN_100; // @[Cat.scala 29:58]
  wire  _GEN_102 = 8'h66 == _T_5[7:0] ? content_102 : _GEN_101; // @[Cat.scala 29:58]
  wire  _GEN_103 = 8'h67 == _T_5[7:0] ? content_103 : _GEN_102; // @[Cat.scala 29:58]
  wire  _GEN_104 = 8'h68 == _T_5[7:0] ? content_104 : _GEN_103; // @[Cat.scala 29:58]
  wire  _GEN_105 = 8'h69 == _T_5[7:0] ? content_105 : _GEN_104; // @[Cat.scala 29:58]
  wire  _GEN_106 = 8'h6a == _T_5[7:0] ? content_106 : _GEN_105; // @[Cat.scala 29:58]
  wire  _GEN_107 = 8'h6b == _T_5[7:0] ? content_107 : _GEN_106; // @[Cat.scala 29:58]
  wire  _GEN_108 = 8'h6c == _T_5[7:0] ? content_108 : _GEN_107; // @[Cat.scala 29:58]
  wire  _GEN_109 = 8'h6d == _T_5[7:0] ? content_109 : _GEN_108; // @[Cat.scala 29:58]
  wire  _GEN_110 = 8'h6e == _T_5[7:0] ? content_110 : _GEN_109; // @[Cat.scala 29:58]
  wire  _GEN_111 = 8'h6f == _T_5[7:0] ? content_111 : _GEN_110; // @[Cat.scala 29:58]
  wire  _GEN_112 = 8'h70 == _T_5[7:0] ? content_112 : _GEN_111; // @[Cat.scala 29:58]
  wire  _GEN_113 = 8'h71 == _T_5[7:0] ? content_113 : _GEN_112; // @[Cat.scala 29:58]
  wire  _GEN_114 = 8'h72 == _T_5[7:0] ? content_114 : _GEN_113; // @[Cat.scala 29:58]
  wire  _GEN_115 = 8'h73 == _T_5[7:0] ? content_115 : _GEN_114; // @[Cat.scala 29:58]
  wire  _GEN_116 = 8'h74 == _T_5[7:0] ? content_116 : _GEN_115; // @[Cat.scala 29:58]
  wire  _GEN_117 = 8'h75 == _T_5[7:0] ? content_117 : _GEN_116; // @[Cat.scala 29:58]
  wire  _GEN_118 = 8'h76 == _T_5[7:0] ? content_118 : _GEN_117; // @[Cat.scala 29:58]
  wire  _GEN_119 = 8'h77 == _T_5[7:0] ? content_119 : _GEN_118; // @[Cat.scala 29:58]
  wire  _GEN_120 = 8'h78 == _T_5[7:0] ? content_120 : _GEN_119; // @[Cat.scala 29:58]
  wire  _GEN_121 = 8'h79 == _T_5[7:0] ? content_121 : _GEN_120; // @[Cat.scala 29:58]
  wire  _GEN_122 = 8'h7a == _T_5[7:0] ? content_122 : _GEN_121; // @[Cat.scala 29:58]
  wire  _GEN_123 = 8'h7b == _T_5[7:0] ? content_123 : _GEN_122; // @[Cat.scala 29:58]
  wire  _GEN_124 = 8'h7c == _T_5[7:0] ? content_124 : _GEN_123; // @[Cat.scala 29:58]
  wire  _GEN_125 = 8'h7d == _T_5[7:0] ? content_125 : _GEN_124; // @[Cat.scala 29:58]
  wire  _GEN_126 = 8'h7e == _T_5[7:0] ? content_126 : _GEN_125; // @[Cat.scala 29:58]
  wire  _GEN_127 = 8'h7f == _T_5[7:0] ? content_127 : _GEN_126; // @[Cat.scala 29:58]
  wire  _GEN_128 = 8'h80 == _T_5[7:0] ? content_128 : _GEN_127; // @[Cat.scala 29:58]
  wire  _GEN_129 = 8'h81 == _T_5[7:0] ? content_129 : _GEN_128; // @[Cat.scala 29:58]
  wire  _GEN_130 = 8'h82 == _T_5[7:0] ? content_130 : _GEN_129; // @[Cat.scala 29:58]
  wire  _GEN_131 = 8'h83 == _T_5[7:0] ? content_131 : _GEN_130; // @[Cat.scala 29:58]
  wire  _GEN_132 = 8'h84 == _T_5[7:0] ? content_132 : _GEN_131; // @[Cat.scala 29:58]
  wire  _GEN_133 = 8'h85 == _T_5[7:0] ? content_133 : _GEN_132; // @[Cat.scala 29:58]
  wire  _GEN_134 = 8'h86 == _T_5[7:0] ? content_134 : _GEN_133; // @[Cat.scala 29:58]
  wire  _GEN_135 = 8'h87 == _T_5[7:0] ? content_135 : _GEN_134; // @[Cat.scala 29:58]
  wire  _GEN_136 = 8'h88 == _T_5[7:0] ? content_136 : _GEN_135; // @[Cat.scala 29:58]
  wire  _GEN_137 = 8'h89 == _T_5[7:0] ? content_137 : _GEN_136; // @[Cat.scala 29:58]
  wire  _GEN_138 = 8'h8a == _T_5[7:0] ? content_138 : _GEN_137; // @[Cat.scala 29:58]
  wire  _GEN_139 = 8'h8b == _T_5[7:0] ? content_139 : _GEN_138; // @[Cat.scala 29:58]
  wire  _GEN_140 = 8'h8c == _T_5[7:0] ? content_140 : _GEN_139; // @[Cat.scala 29:58]
  wire  _GEN_141 = 8'h8d == _T_5[7:0] ? content_141 : _GEN_140; // @[Cat.scala 29:58]
  wire  _GEN_142 = 8'h8e == _T_5[7:0] ? content_142 : _GEN_141; // @[Cat.scala 29:58]
  wire  _GEN_143 = 8'h8f == _T_5[7:0] ? content_143 : _GEN_142; // @[Cat.scala 29:58]
  wire  _GEN_144 = 8'h90 == _T_5[7:0] ? content_144 : _GEN_143; // @[Cat.scala 29:58]
  wire  _GEN_145 = 8'h91 == _T_5[7:0] ? content_145 : _GEN_144; // @[Cat.scala 29:58]
  wire  _GEN_146 = 8'h92 == _T_5[7:0] ? content_146 : _GEN_145; // @[Cat.scala 29:58]
  wire  _GEN_147 = 8'h93 == _T_5[7:0] ? content_147 : _GEN_146; // @[Cat.scala 29:58]
  wire  _GEN_148 = 8'h94 == _T_5[7:0] ? content_148 : _GEN_147; // @[Cat.scala 29:58]
  wire  _GEN_149 = 8'h95 == _T_5[7:0] ? content_149 : _GEN_148; // @[Cat.scala 29:58]
  wire  _GEN_150 = 8'h96 == _T_5[7:0] ? content_150 : _GEN_149; // @[Cat.scala 29:58]
  wire  _GEN_151 = 8'h97 == _T_5[7:0] ? content_151 : _GEN_150; // @[Cat.scala 29:58]
  wire  _GEN_152 = 8'h98 == _T_5[7:0] ? content_152 : _GEN_151; // @[Cat.scala 29:58]
  wire  _GEN_153 = 8'h99 == _T_5[7:0] ? content_153 : _GEN_152; // @[Cat.scala 29:58]
  wire  _GEN_154 = 8'h9a == _T_5[7:0] ? content_154 : _GEN_153; // @[Cat.scala 29:58]
  wire  _GEN_155 = 8'h9b == _T_5[7:0] ? content_155 : _GEN_154; // @[Cat.scala 29:58]
  wire  _GEN_156 = 8'h9c == _T_5[7:0] ? content_156 : _GEN_155; // @[Cat.scala 29:58]
  wire  _GEN_157 = 8'h9d == _T_5[7:0] ? content_157 : _GEN_156; // @[Cat.scala 29:58]
  wire  _GEN_158 = 8'h9e == _T_5[7:0] ? content_158 : _GEN_157; // @[Cat.scala 29:58]
  wire  _GEN_159 = 8'h9f == _T_5[7:0] ? content_159 : _GEN_158; // @[Cat.scala 29:58]
  wire  _GEN_160 = 8'ha0 == _T_5[7:0] ? content_160 : _GEN_159; // @[Cat.scala 29:58]
  wire  _GEN_161 = 8'ha1 == _T_5[7:0] ? content_161 : _GEN_160; // @[Cat.scala 29:58]
  wire  _GEN_162 = 8'ha2 == _T_5[7:0] ? content_162 : _GEN_161; // @[Cat.scala 29:58]
  wire  _GEN_163 = 8'ha3 == _T_5[7:0] ? content_163 : _GEN_162; // @[Cat.scala 29:58]
  wire  _GEN_164 = 8'ha4 == _T_5[7:0] ? content_164 : _GEN_163; // @[Cat.scala 29:58]
  wire  _GEN_165 = 8'ha5 == _T_5[7:0] ? content_165 : _GEN_164; // @[Cat.scala 29:58]
  wire  _GEN_166 = 8'ha6 == _T_5[7:0] ? content_166 : _GEN_165; // @[Cat.scala 29:58]
  wire  _GEN_167 = 8'ha7 == _T_5[7:0] ? content_167 : _GEN_166; // @[Cat.scala 29:58]
  wire  _GEN_168 = 8'ha8 == _T_5[7:0] ? content_168 : _GEN_167; // @[Cat.scala 29:58]
  wire  _GEN_169 = 8'ha9 == _T_5[7:0] ? content_169 : _GEN_168; // @[Cat.scala 29:58]
  wire  _GEN_170 = 8'haa == _T_5[7:0] ? content_170 : _GEN_169; // @[Cat.scala 29:58]
  wire  _GEN_171 = 8'hab == _T_5[7:0] ? content_171 : _GEN_170; // @[Cat.scala 29:58]
  wire  _GEN_172 = 8'hac == _T_5[7:0] ? content_172 : _GEN_171; // @[Cat.scala 29:58]
  wire  _GEN_173 = 8'had == _T_5[7:0] ? content_173 : _GEN_172; // @[Cat.scala 29:58]
  wire  _GEN_174 = 8'hae == _T_5[7:0] ? content_174 : _GEN_173; // @[Cat.scala 29:58]
  wire  _GEN_175 = 8'haf == _T_5[7:0] ? content_175 : _GEN_174; // @[Cat.scala 29:58]
  wire  _GEN_176 = 8'hb0 == _T_5[7:0] ? content_176 : _GEN_175; // @[Cat.scala 29:58]
  wire  _GEN_177 = 8'hb1 == _T_5[7:0] ? content_177 : _GEN_176; // @[Cat.scala 29:58]
  wire  _GEN_178 = 8'hb2 == _T_5[7:0] ? content_178 : _GEN_177; // @[Cat.scala 29:58]
  wire  _GEN_179 = 8'hb3 == _T_5[7:0] ? content_179 : _GEN_178; // @[Cat.scala 29:58]
  wire  _GEN_180 = 8'hb4 == _T_5[7:0] ? content_180 : _GEN_179; // @[Cat.scala 29:58]
  wire  _GEN_181 = 8'hb5 == _T_5[7:0] ? content_181 : _GEN_180; // @[Cat.scala 29:58]
  wire  _GEN_182 = 8'hb6 == _T_5[7:0] ? content_182 : _GEN_181; // @[Cat.scala 29:58]
  wire  _GEN_183 = 8'hb7 == _T_5[7:0] ? content_183 : _GEN_182; // @[Cat.scala 29:58]
  wire  _GEN_184 = 8'hb8 == _T_5[7:0] ? content_184 : _GEN_183; // @[Cat.scala 29:58]
  wire  _GEN_185 = 8'hb9 == _T_5[7:0] ? content_185 : _GEN_184; // @[Cat.scala 29:58]
  wire  _GEN_186 = 8'hba == _T_5[7:0] ? content_186 : _GEN_185; // @[Cat.scala 29:58]
  wire  _GEN_187 = 8'hbb == _T_5[7:0] ? content_187 : _GEN_186; // @[Cat.scala 29:58]
  wire  _GEN_188 = 8'hbc == _T_5[7:0] ? content_188 : _GEN_187; // @[Cat.scala 29:58]
  wire  _GEN_189 = 8'hbd == _T_5[7:0] ? content_189 : _GEN_188; // @[Cat.scala 29:58]
  wire  _GEN_190 = 8'hbe == _T_5[7:0] ? content_190 : _GEN_189; // @[Cat.scala 29:58]
  wire  _GEN_191 = 8'hbf == _T_5[7:0] ? content_191 : _GEN_190; // @[Cat.scala 29:58]
  wire  _GEN_192 = 8'hc0 == _T_5[7:0] ? content_192 : _GEN_191; // @[Cat.scala 29:58]
  wire  _GEN_193 = 8'hc1 == _T_5[7:0] ? content_193 : _GEN_192; // @[Cat.scala 29:58]
  wire  _GEN_194 = 8'hc2 == _T_5[7:0] ? content_194 : _GEN_193; // @[Cat.scala 29:58]
  wire  _GEN_195 = 8'hc3 == _T_5[7:0] ? content_195 : _GEN_194; // @[Cat.scala 29:58]
  wire  _GEN_196 = 8'hc4 == _T_5[7:0] ? content_196 : _GEN_195; // @[Cat.scala 29:58]
  wire  _GEN_197 = 8'hc5 == _T_5[7:0] ? content_197 : _GEN_196; // @[Cat.scala 29:58]
  wire  _GEN_198 = 8'hc6 == _T_5[7:0] ? content_198 : _GEN_197; // @[Cat.scala 29:58]
  wire  _GEN_199 = 8'hc7 == _T_5[7:0] ? content_199 : _GEN_198; // @[Cat.scala 29:58]
  wire  _GEN_200 = 8'hc8 == _T_5[7:0] ? content_200 : _GEN_199; // @[Cat.scala 29:58]
  wire  _GEN_201 = 8'hc9 == _T_5[7:0] ? content_201 : _GEN_200; // @[Cat.scala 29:58]
  wire  _GEN_202 = 8'hca == _T_5[7:0] ? content_202 : _GEN_201; // @[Cat.scala 29:58]
  wire  _GEN_203 = 8'hcb == _T_5[7:0] ? content_203 : _GEN_202; // @[Cat.scala 29:58]
  wire  _GEN_204 = 8'hcc == _T_5[7:0] ? content_204 : _GEN_203; // @[Cat.scala 29:58]
  wire  _GEN_205 = 8'hcd == _T_5[7:0] ? content_205 : _GEN_204; // @[Cat.scala 29:58]
  wire  _GEN_206 = 8'hce == _T_5[7:0] ? content_206 : _GEN_205; // @[Cat.scala 29:58]
  wire  _GEN_207 = 8'hcf == _T_5[7:0] ? content_207 : _GEN_206; // @[Cat.scala 29:58]
  wire  _GEN_208 = 8'hd0 == _T_5[7:0] ? content_208 : _GEN_207; // @[Cat.scala 29:58]
  wire  _GEN_209 = 8'hd1 == _T_5[7:0] ? content_209 : _GEN_208; // @[Cat.scala 29:58]
  wire  _GEN_210 = 8'hd2 == _T_5[7:0] ? content_210 : _GEN_209; // @[Cat.scala 29:58]
  wire  _GEN_211 = 8'hd3 == _T_5[7:0] ? content_211 : _GEN_210; // @[Cat.scala 29:58]
  wire  _GEN_212 = 8'hd4 == _T_5[7:0] ? content_212 : _GEN_211; // @[Cat.scala 29:58]
  wire  _GEN_213 = 8'hd5 == _T_5[7:0] ? content_213 : _GEN_212; // @[Cat.scala 29:58]
  wire  _GEN_214 = 8'hd6 == _T_5[7:0] ? content_214 : _GEN_213; // @[Cat.scala 29:58]
  wire  _GEN_215 = 8'hd7 == _T_5[7:0] ? content_215 : _GEN_214; // @[Cat.scala 29:58]
  wire  _GEN_216 = 8'hd8 == _T_5[7:0] ? content_216 : _GEN_215; // @[Cat.scala 29:58]
  wire  _GEN_217 = 8'hd9 == _T_5[7:0] ? content_217 : _GEN_216; // @[Cat.scala 29:58]
  wire  _GEN_218 = 8'hda == _T_5[7:0] ? content_218 : _GEN_217; // @[Cat.scala 29:58]
  wire  _GEN_219 = 8'hdb == _T_5[7:0] ? content_219 : _GEN_218; // @[Cat.scala 29:58]
  wire  _GEN_220 = 8'hdc == _T_5[7:0] ? content_220 : _GEN_219; // @[Cat.scala 29:58]
  wire  _GEN_221 = 8'hdd == _T_5[7:0] ? content_221 : _GEN_220; // @[Cat.scala 29:58]
  wire  _GEN_222 = 8'hde == _T_5[7:0] ? content_222 : _GEN_221; // @[Cat.scala 29:58]
  wire  _GEN_223 = 8'hdf == _T_5[7:0] ? content_223 : _GEN_222; // @[Cat.scala 29:58]
  wire  _GEN_224 = 8'he0 == _T_5[7:0] ? content_224 : _GEN_223; // @[Cat.scala 29:58]
  wire  _GEN_225 = 8'he1 == _T_5[7:0] ? content_225 : _GEN_224; // @[Cat.scala 29:58]
  wire  _GEN_226 = 8'he2 == _T_5[7:0] ? content_226 : _GEN_225; // @[Cat.scala 29:58]
  wire  _GEN_227 = 8'he3 == _T_5[7:0] ? content_227 : _GEN_226; // @[Cat.scala 29:58]
  wire  _GEN_228 = 8'he4 == _T_5[7:0] ? content_228 : _GEN_227; // @[Cat.scala 29:58]
  wire  _GEN_229 = 8'he5 == _T_5[7:0] ? content_229 : _GEN_228; // @[Cat.scala 29:58]
  wire  _GEN_230 = 8'he6 == _T_5[7:0] ? content_230 : _GEN_229; // @[Cat.scala 29:58]
  wire  _GEN_231 = 8'he7 == _T_5[7:0] ? content_231 : _GEN_230; // @[Cat.scala 29:58]
  wire  _GEN_232 = 8'he8 == _T_5[7:0] ? content_232 : _GEN_231; // @[Cat.scala 29:58]
  wire  _GEN_233 = 8'he9 == _T_5[7:0] ? content_233 : _GEN_232; // @[Cat.scala 29:58]
  wire  _GEN_234 = 8'hea == _T_5[7:0] ? content_234 : _GEN_233; // @[Cat.scala 29:58]
  wire  _GEN_235 = 8'heb == _T_5[7:0] ? content_235 : _GEN_234; // @[Cat.scala 29:58]
  wire  _GEN_236 = 8'hec == _T_5[7:0] ? content_236 : _GEN_235; // @[Cat.scala 29:58]
  wire  _GEN_237 = 8'hed == _T_5[7:0] ? content_237 : _GEN_236; // @[Cat.scala 29:58]
  wire  _GEN_238 = 8'hee == _T_5[7:0] ? content_238 : _GEN_237; // @[Cat.scala 29:58]
  wire  _GEN_239 = 8'hef == _T_5[7:0] ? content_239 : _GEN_238; // @[Cat.scala 29:58]
  wire  _GEN_240 = 8'hf0 == _T_5[7:0] ? content_240 : _GEN_239; // @[Cat.scala 29:58]
  wire  _GEN_241 = 8'hf1 == _T_5[7:0] ? content_241 : _GEN_240; // @[Cat.scala 29:58]
  wire  _GEN_242 = 8'hf2 == _T_5[7:0] ? content_242 : _GEN_241; // @[Cat.scala 29:58]
  wire  _GEN_243 = 8'hf3 == _T_5[7:0] ? content_243 : _GEN_242; // @[Cat.scala 29:58]
  wire  _GEN_244 = 8'hf4 == _T_5[7:0] ? content_244 : _GEN_243; // @[Cat.scala 29:58]
  wire  _GEN_245 = 8'hf5 == _T_5[7:0] ? content_245 : _GEN_244; // @[Cat.scala 29:58]
  wire  _GEN_246 = 8'hf6 == _T_5[7:0] ? content_246 : _GEN_245; // @[Cat.scala 29:58]
  wire  _GEN_247 = 8'hf7 == _T_5[7:0] ? content_247 : _GEN_246; // @[Cat.scala 29:58]
  wire  _GEN_248 = 8'hf8 == _T_5[7:0] ? content_248 : _GEN_247; // @[Cat.scala 29:58]
  wire  _GEN_249 = 8'hf9 == _T_5[7:0] ? content_249 : _GEN_248; // @[Cat.scala 29:58]
  wire  _GEN_250 = 8'hfa == _T_5[7:0] ? content_250 : _GEN_249; // @[Cat.scala 29:58]
  wire  _GEN_251 = 8'hfb == _T_5[7:0] ? content_251 : _GEN_250; // @[Cat.scala 29:58]
  wire  _GEN_252 = 8'hfc == _T_5[7:0] ? content_252 : _GEN_251; // @[Cat.scala 29:58]
  wire  _GEN_253 = 8'hfd == _T_5[7:0] ? content_253 : _GEN_252; // @[Cat.scala 29:58]
  wire  _GEN_254 = 8'hfe == _T_5[7:0] ? content_254 : _GEN_253; // @[Cat.scala 29:58]
  wire  _GEN_255 = 8'hff == _T_5[7:0] ? content_255 : _GEN_254; // @[Cat.scala 29:58]
  wire  _GEN_257 = 8'h1 == _T_1[7:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_258 = 8'h2 == _T_1[7:0] ? content_2 : _GEN_257; // @[Cat.scala 29:58]
  wire  _GEN_259 = 8'h3 == _T_1[7:0] ? content_3 : _GEN_258; // @[Cat.scala 29:58]
  wire  _GEN_260 = 8'h4 == _T_1[7:0] ? content_4 : _GEN_259; // @[Cat.scala 29:58]
  wire  _GEN_261 = 8'h5 == _T_1[7:0] ? content_5 : _GEN_260; // @[Cat.scala 29:58]
  wire  _GEN_262 = 8'h6 == _T_1[7:0] ? content_6 : _GEN_261; // @[Cat.scala 29:58]
  wire  _GEN_263 = 8'h7 == _T_1[7:0] ? content_7 : _GEN_262; // @[Cat.scala 29:58]
  wire  _GEN_264 = 8'h8 == _T_1[7:0] ? content_8 : _GEN_263; // @[Cat.scala 29:58]
  wire  _GEN_265 = 8'h9 == _T_1[7:0] ? content_9 : _GEN_264; // @[Cat.scala 29:58]
  wire  _GEN_266 = 8'ha == _T_1[7:0] ? content_10 : _GEN_265; // @[Cat.scala 29:58]
  wire  _GEN_267 = 8'hb == _T_1[7:0] ? content_11 : _GEN_266; // @[Cat.scala 29:58]
  wire  _GEN_268 = 8'hc == _T_1[7:0] ? content_12 : _GEN_267; // @[Cat.scala 29:58]
  wire  _GEN_269 = 8'hd == _T_1[7:0] ? content_13 : _GEN_268; // @[Cat.scala 29:58]
  wire  _GEN_270 = 8'he == _T_1[7:0] ? content_14 : _GEN_269; // @[Cat.scala 29:58]
  wire  _GEN_271 = 8'hf == _T_1[7:0] ? content_15 : _GEN_270; // @[Cat.scala 29:58]
  wire  _GEN_272 = 8'h10 == _T_1[7:0] ? content_16 : _GEN_271; // @[Cat.scala 29:58]
  wire  _GEN_273 = 8'h11 == _T_1[7:0] ? content_17 : _GEN_272; // @[Cat.scala 29:58]
  wire  _GEN_274 = 8'h12 == _T_1[7:0] ? content_18 : _GEN_273; // @[Cat.scala 29:58]
  wire  _GEN_275 = 8'h13 == _T_1[7:0] ? content_19 : _GEN_274; // @[Cat.scala 29:58]
  wire  _GEN_276 = 8'h14 == _T_1[7:0] ? content_20 : _GEN_275; // @[Cat.scala 29:58]
  wire  _GEN_277 = 8'h15 == _T_1[7:0] ? content_21 : _GEN_276; // @[Cat.scala 29:58]
  wire  _GEN_278 = 8'h16 == _T_1[7:0] ? content_22 : _GEN_277; // @[Cat.scala 29:58]
  wire  _GEN_279 = 8'h17 == _T_1[7:0] ? content_23 : _GEN_278; // @[Cat.scala 29:58]
  wire  _GEN_280 = 8'h18 == _T_1[7:0] ? content_24 : _GEN_279; // @[Cat.scala 29:58]
  wire  _GEN_281 = 8'h19 == _T_1[7:0] ? content_25 : _GEN_280; // @[Cat.scala 29:58]
  wire  _GEN_282 = 8'h1a == _T_1[7:0] ? content_26 : _GEN_281; // @[Cat.scala 29:58]
  wire  _GEN_283 = 8'h1b == _T_1[7:0] ? content_27 : _GEN_282; // @[Cat.scala 29:58]
  wire  _GEN_284 = 8'h1c == _T_1[7:0] ? content_28 : _GEN_283; // @[Cat.scala 29:58]
  wire  _GEN_285 = 8'h1d == _T_1[7:0] ? content_29 : _GEN_284; // @[Cat.scala 29:58]
  wire  _GEN_286 = 8'h1e == _T_1[7:0] ? content_30 : _GEN_285; // @[Cat.scala 29:58]
  wire  _GEN_287 = 8'h1f == _T_1[7:0] ? content_31 : _GEN_286; // @[Cat.scala 29:58]
  wire  _GEN_288 = 8'h20 == _T_1[7:0] ? content_32 : _GEN_287; // @[Cat.scala 29:58]
  wire  _GEN_289 = 8'h21 == _T_1[7:0] ? content_33 : _GEN_288; // @[Cat.scala 29:58]
  wire  _GEN_290 = 8'h22 == _T_1[7:0] ? content_34 : _GEN_289; // @[Cat.scala 29:58]
  wire  _GEN_291 = 8'h23 == _T_1[7:0] ? content_35 : _GEN_290; // @[Cat.scala 29:58]
  wire  _GEN_292 = 8'h24 == _T_1[7:0] ? content_36 : _GEN_291; // @[Cat.scala 29:58]
  wire  _GEN_293 = 8'h25 == _T_1[7:0] ? content_37 : _GEN_292; // @[Cat.scala 29:58]
  wire  _GEN_294 = 8'h26 == _T_1[7:0] ? content_38 : _GEN_293; // @[Cat.scala 29:58]
  wire  _GEN_295 = 8'h27 == _T_1[7:0] ? content_39 : _GEN_294; // @[Cat.scala 29:58]
  wire  _GEN_296 = 8'h28 == _T_1[7:0] ? content_40 : _GEN_295; // @[Cat.scala 29:58]
  wire  _GEN_297 = 8'h29 == _T_1[7:0] ? content_41 : _GEN_296; // @[Cat.scala 29:58]
  wire  _GEN_298 = 8'h2a == _T_1[7:0] ? content_42 : _GEN_297; // @[Cat.scala 29:58]
  wire  _GEN_299 = 8'h2b == _T_1[7:0] ? content_43 : _GEN_298; // @[Cat.scala 29:58]
  wire  _GEN_300 = 8'h2c == _T_1[7:0] ? content_44 : _GEN_299; // @[Cat.scala 29:58]
  wire  _GEN_301 = 8'h2d == _T_1[7:0] ? content_45 : _GEN_300; // @[Cat.scala 29:58]
  wire  _GEN_302 = 8'h2e == _T_1[7:0] ? content_46 : _GEN_301; // @[Cat.scala 29:58]
  wire  _GEN_303 = 8'h2f == _T_1[7:0] ? content_47 : _GEN_302; // @[Cat.scala 29:58]
  wire  _GEN_304 = 8'h30 == _T_1[7:0] ? content_48 : _GEN_303; // @[Cat.scala 29:58]
  wire  _GEN_305 = 8'h31 == _T_1[7:0] ? content_49 : _GEN_304; // @[Cat.scala 29:58]
  wire  _GEN_306 = 8'h32 == _T_1[7:0] ? content_50 : _GEN_305; // @[Cat.scala 29:58]
  wire  _GEN_307 = 8'h33 == _T_1[7:0] ? content_51 : _GEN_306; // @[Cat.scala 29:58]
  wire  _GEN_308 = 8'h34 == _T_1[7:0] ? content_52 : _GEN_307; // @[Cat.scala 29:58]
  wire  _GEN_309 = 8'h35 == _T_1[7:0] ? content_53 : _GEN_308; // @[Cat.scala 29:58]
  wire  _GEN_310 = 8'h36 == _T_1[7:0] ? content_54 : _GEN_309; // @[Cat.scala 29:58]
  wire  _GEN_311 = 8'h37 == _T_1[7:0] ? content_55 : _GEN_310; // @[Cat.scala 29:58]
  wire  _GEN_312 = 8'h38 == _T_1[7:0] ? content_56 : _GEN_311; // @[Cat.scala 29:58]
  wire  _GEN_313 = 8'h39 == _T_1[7:0] ? content_57 : _GEN_312; // @[Cat.scala 29:58]
  wire  _GEN_314 = 8'h3a == _T_1[7:0] ? content_58 : _GEN_313; // @[Cat.scala 29:58]
  wire  _GEN_315 = 8'h3b == _T_1[7:0] ? content_59 : _GEN_314; // @[Cat.scala 29:58]
  wire  _GEN_316 = 8'h3c == _T_1[7:0] ? content_60 : _GEN_315; // @[Cat.scala 29:58]
  wire  _GEN_317 = 8'h3d == _T_1[7:0] ? content_61 : _GEN_316; // @[Cat.scala 29:58]
  wire  _GEN_318 = 8'h3e == _T_1[7:0] ? content_62 : _GEN_317; // @[Cat.scala 29:58]
  wire  _GEN_319 = 8'h3f == _T_1[7:0] ? content_63 : _GEN_318; // @[Cat.scala 29:58]
  wire  _GEN_320 = 8'h40 == _T_1[7:0] ? content_64 : _GEN_319; // @[Cat.scala 29:58]
  wire  _GEN_321 = 8'h41 == _T_1[7:0] ? content_65 : _GEN_320; // @[Cat.scala 29:58]
  wire  _GEN_322 = 8'h42 == _T_1[7:0] ? content_66 : _GEN_321; // @[Cat.scala 29:58]
  wire  _GEN_323 = 8'h43 == _T_1[7:0] ? content_67 : _GEN_322; // @[Cat.scala 29:58]
  wire  _GEN_324 = 8'h44 == _T_1[7:0] ? content_68 : _GEN_323; // @[Cat.scala 29:58]
  wire  _GEN_325 = 8'h45 == _T_1[7:0] ? content_69 : _GEN_324; // @[Cat.scala 29:58]
  wire  _GEN_326 = 8'h46 == _T_1[7:0] ? content_70 : _GEN_325; // @[Cat.scala 29:58]
  wire  _GEN_327 = 8'h47 == _T_1[7:0] ? content_71 : _GEN_326; // @[Cat.scala 29:58]
  wire  _GEN_328 = 8'h48 == _T_1[7:0] ? content_72 : _GEN_327; // @[Cat.scala 29:58]
  wire  _GEN_329 = 8'h49 == _T_1[7:0] ? content_73 : _GEN_328; // @[Cat.scala 29:58]
  wire  _GEN_330 = 8'h4a == _T_1[7:0] ? content_74 : _GEN_329; // @[Cat.scala 29:58]
  wire  _GEN_331 = 8'h4b == _T_1[7:0] ? content_75 : _GEN_330; // @[Cat.scala 29:58]
  wire  _GEN_332 = 8'h4c == _T_1[7:0] ? content_76 : _GEN_331; // @[Cat.scala 29:58]
  wire  _GEN_333 = 8'h4d == _T_1[7:0] ? content_77 : _GEN_332; // @[Cat.scala 29:58]
  wire  _GEN_334 = 8'h4e == _T_1[7:0] ? content_78 : _GEN_333; // @[Cat.scala 29:58]
  wire  _GEN_335 = 8'h4f == _T_1[7:0] ? content_79 : _GEN_334; // @[Cat.scala 29:58]
  wire  _GEN_336 = 8'h50 == _T_1[7:0] ? content_80 : _GEN_335; // @[Cat.scala 29:58]
  wire  _GEN_337 = 8'h51 == _T_1[7:0] ? content_81 : _GEN_336; // @[Cat.scala 29:58]
  wire  _GEN_338 = 8'h52 == _T_1[7:0] ? content_82 : _GEN_337; // @[Cat.scala 29:58]
  wire  _GEN_339 = 8'h53 == _T_1[7:0] ? content_83 : _GEN_338; // @[Cat.scala 29:58]
  wire  _GEN_340 = 8'h54 == _T_1[7:0] ? content_84 : _GEN_339; // @[Cat.scala 29:58]
  wire  _GEN_341 = 8'h55 == _T_1[7:0] ? content_85 : _GEN_340; // @[Cat.scala 29:58]
  wire  _GEN_342 = 8'h56 == _T_1[7:0] ? content_86 : _GEN_341; // @[Cat.scala 29:58]
  wire  _GEN_343 = 8'h57 == _T_1[7:0] ? content_87 : _GEN_342; // @[Cat.scala 29:58]
  wire  _GEN_344 = 8'h58 == _T_1[7:0] ? content_88 : _GEN_343; // @[Cat.scala 29:58]
  wire  _GEN_345 = 8'h59 == _T_1[7:0] ? content_89 : _GEN_344; // @[Cat.scala 29:58]
  wire  _GEN_346 = 8'h5a == _T_1[7:0] ? content_90 : _GEN_345; // @[Cat.scala 29:58]
  wire  _GEN_347 = 8'h5b == _T_1[7:0] ? content_91 : _GEN_346; // @[Cat.scala 29:58]
  wire  _GEN_348 = 8'h5c == _T_1[7:0] ? content_92 : _GEN_347; // @[Cat.scala 29:58]
  wire  _GEN_349 = 8'h5d == _T_1[7:0] ? content_93 : _GEN_348; // @[Cat.scala 29:58]
  wire  _GEN_350 = 8'h5e == _T_1[7:0] ? content_94 : _GEN_349; // @[Cat.scala 29:58]
  wire  _GEN_351 = 8'h5f == _T_1[7:0] ? content_95 : _GEN_350; // @[Cat.scala 29:58]
  wire  _GEN_352 = 8'h60 == _T_1[7:0] ? content_96 : _GEN_351; // @[Cat.scala 29:58]
  wire  _GEN_353 = 8'h61 == _T_1[7:0] ? content_97 : _GEN_352; // @[Cat.scala 29:58]
  wire  _GEN_354 = 8'h62 == _T_1[7:0] ? content_98 : _GEN_353; // @[Cat.scala 29:58]
  wire  _GEN_355 = 8'h63 == _T_1[7:0] ? content_99 : _GEN_354; // @[Cat.scala 29:58]
  wire  _GEN_356 = 8'h64 == _T_1[7:0] ? content_100 : _GEN_355; // @[Cat.scala 29:58]
  wire  _GEN_357 = 8'h65 == _T_1[7:0] ? content_101 : _GEN_356; // @[Cat.scala 29:58]
  wire  _GEN_358 = 8'h66 == _T_1[7:0] ? content_102 : _GEN_357; // @[Cat.scala 29:58]
  wire  _GEN_359 = 8'h67 == _T_1[7:0] ? content_103 : _GEN_358; // @[Cat.scala 29:58]
  wire  _GEN_360 = 8'h68 == _T_1[7:0] ? content_104 : _GEN_359; // @[Cat.scala 29:58]
  wire  _GEN_361 = 8'h69 == _T_1[7:0] ? content_105 : _GEN_360; // @[Cat.scala 29:58]
  wire  _GEN_362 = 8'h6a == _T_1[7:0] ? content_106 : _GEN_361; // @[Cat.scala 29:58]
  wire  _GEN_363 = 8'h6b == _T_1[7:0] ? content_107 : _GEN_362; // @[Cat.scala 29:58]
  wire  _GEN_364 = 8'h6c == _T_1[7:0] ? content_108 : _GEN_363; // @[Cat.scala 29:58]
  wire  _GEN_365 = 8'h6d == _T_1[7:0] ? content_109 : _GEN_364; // @[Cat.scala 29:58]
  wire  _GEN_366 = 8'h6e == _T_1[7:0] ? content_110 : _GEN_365; // @[Cat.scala 29:58]
  wire  _GEN_367 = 8'h6f == _T_1[7:0] ? content_111 : _GEN_366; // @[Cat.scala 29:58]
  wire  _GEN_368 = 8'h70 == _T_1[7:0] ? content_112 : _GEN_367; // @[Cat.scala 29:58]
  wire  _GEN_369 = 8'h71 == _T_1[7:0] ? content_113 : _GEN_368; // @[Cat.scala 29:58]
  wire  _GEN_370 = 8'h72 == _T_1[7:0] ? content_114 : _GEN_369; // @[Cat.scala 29:58]
  wire  _GEN_371 = 8'h73 == _T_1[7:0] ? content_115 : _GEN_370; // @[Cat.scala 29:58]
  wire  _GEN_372 = 8'h74 == _T_1[7:0] ? content_116 : _GEN_371; // @[Cat.scala 29:58]
  wire  _GEN_373 = 8'h75 == _T_1[7:0] ? content_117 : _GEN_372; // @[Cat.scala 29:58]
  wire  _GEN_374 = 8'h76 == _T_1[7:0] ? content_118 : _GEN_373; // @[Cat.scala 29:58]
  wire  _GEN_375 = 8'h77 == _T_1[7:0] ? content_119 : _GEN_374; // @[Cat.scala 29:58]
  wire  _GEN_376 = 8'h78 == _T_1[7:0] ? content_120 : _GEN_375; // @[Cat.scala 29:58]
  wire  _GEN_377 = 8'h79 == _T_1[7:0] ? content_121 : _GEN_376; // @[Cat.scala 29:58]
  wire  _GEN_378 = 8'h7a == _T_1[7:0] ? content_122 : _GEN_377; // @[Cat.scala 29:58]
  wire  _GEN_379 = 8'h7b == _T_1[7:0] ? content_123 : _GEN_378; // @[Cat.scala 29:58]
  wire  _GEN_380 = 8'h7c == _T_1[7:0] ? content_124 : _GEN_379; // @[Cat.scala 29:58]
  wire  _GEN_381 = 8'h7d == _T_1[7:0] ? content_125 : _GEN_380; // @[Cat.scala 29:58]
  wire  _GEN_382 = 8'h7e == _T_1[7:0] ? content_126 : _GEN_381; // @[Cat.scala 29:58]
  wire  _GEN_383 = 8'h7f == _T_1[7:0] ? content_127 : _GEN_382; // @[Cat.scala 29:58]
  wire  _GEN_384 = 8'h80 == _T_1[7:0] ? content_128 : _GEN_383; // @[Cat.scala 29:58]
  wire  _GEN_385 = 8'h81 == _T_1[7:0] ? content_129 : _GEN_384; // @[Cat.scala 29:58]
  wire  _GEN_386 = 8'h82 == _T_1[7:0] ? content_130 : _GEN_385; // @[Cat.scala 29:58]
  wire  _GEN_387 = 8'h83 == _T_1[7:0] ? content_131 : _GEN_386; // @[Cat.scala 29:58]
  wire  _GEN_388 = 8'h84 == _T_1[7:0] ? content_132 : _GEN_387; // @[Cat.scala 29:58]
  wire  _GEN_389 = 8'h85 == _T_1[7:0] ? content_133 : _GEN_388; // @[Cat.scala 29:58]
  wire  _GEN_390 = 8'h86 == _T_1[7:0] ? content_134 : _GEN_389; // @[Cat.scala 29:58]
  wire  _GEN_391 = 8'h87 == _T_1[7:0] ? content_135 : _GEN_390; // @[Cat.scala 29:58]
  wire  _GEN_392 = 8'h88 == _T_1[7:0] ? content_136 : _GEN_391; // @[Cat.scala 29:58]
  wire  _GEN_393 = 8'h89 == _T_1[7:0] ? content_137 : _GEN_392; // @[Cat.scala 29:58]
  wire  _GEN_394 = 8'h8a == _T_1[7:0] ? content_138 : _GEN_393; // @[Cat.scala 29:58]
  wire  _GEN_395 = 8'h8b == _T_1[7:0] ? content_139 : _GEN_394; // @[Cat.scala 29:58]
  wire  _GEN_396 = 8'h8c == _T_1[7:0] ? content_140 : _GEN_395; // @[Cat.scala 29:58]
  wire  _GEN_397 = 8'h8d == _T_1[7:0] ? content_141 : _GEN_396; // @[Cat.scala 29:58]
  wire  _GEN_398 = 8'h8e == _T_1[7:0] ? content_142 : _GEN_397; // @[Cat.scala 29:58]
  wire  _GEN_399 = 8'h8f == _T_1[7:0] ? content_143 : _GEN_398; // @[Cat.scala 29:58]
  wire  _GEN_400 = 8'h90 == _T_1[7:0] ? content_144 : _GEN_399; // @[Cat.scala 29:58]
  wire  _GEN_401 = 8'h91 == _T_1[7:0] ? content_145 : _GEN_400; // @[Cat.scala 29:58]
  wire  _GEN_402 = 8'h92 == _T_1[7:0] ? content_146 : _GEN_401; // @[Cat.scala 29:58]
  wire  _GEN_403 = 8'h93 == _T_1[7:0] ? content_147 : _GEN_402; // @[Cat.scala 29:58]
  wire  _GEN_404 = 8'h94 == _T_1[7:0] ? content_148 : _GEN_403; // @[Cat.scala 29:58]
  wire  _GEN_405 = 8'h95 == _T_1[7:0] ? content_149 : _GEN_404; // @[Cat.scala 29:58]
  wire  _GEN_406 = 8'h96 == _T_1[7:0] ? content_150 : _GEN_405; // @[Cat.scala 29:58]
  wire  _GEN_407 = 8'h97 == _T_1[7:0] ? content_151 : _GEN_406; // @[Cat.scala 29:58]
  wire  _GEN_408 = 8'h98 == _T_1[7:0] ? content_152 : _GEN_407; // @[Cat.scala 29:58]
  wire  _GEN_409 = 8'h99 == _T_1[7:0] ? content_153 : _GEN_408; // @[Cat.scala 29:58]
  wire  _GEN_410 = 8'h9a == _T_1[7:0] ? content_154 : _GEN_409; // @[Cat.scala 29:58]
  wire  _GEN_411 = 8'h9b == _T_1[7:0] ? content_155 : _GEN_410; // @[Cat.scala 29:58]
  wire  _GEN_412 = 8'h9c == _T_1[7:0] ? content_156 : _GEN_411; // @[Cat.scala 29:58]
  wire  _GEN_413 = 8'h9d == _T_1[7:0] ? content_157 : _GEN_412; // @[Cat.scala 29:58]
  wire  _GEN_414 = 8'h9e == _T_1[7:0] ? content_158 : _GEN_413; // @[Cat.scala 29:58]
  wire  _GEN_415 = 8'h9f == _T_1[7:0] ? content_159 : _GEN_414; // @[Cat.scala 29:58]
  wire  _GEN_416 = 8'ha0 == _T_1[7:0] ? content_160 : _GEN_415; // @[Cat.scala 29:58]
  wire  _GEN_417 = 8'ha1 == _T_1[7:0] ? content_161 : _GEN_416; // @[Cat.scala 29:58]
  wire  _GEN_418 = 8'ha2 == _T_1[7:0] ? content_162 : _GEN_417; // @[Cat.scala 29:58]
  wire  _GEN_419 = 8'ha3 == _T_1[7:0] ? content_163 : _GEN_418; // @[Cat.scala 29:58]
  wire  _GEN_420 = 8'ha4 == _T_1[7:0] ? content_164 : _GEN_419; // @[Cat.scala 29:58]
  wire  _GEN_421 = 8'ha5 == _T_1[7:0] ? content_165 : _GEN_420; // @[Cat.scala 29:58]
  wire  _GEN_422 = 8'ha6 == _T_1[7:0] ? content_166 : _GEN_421; // @[Cat.scala 29:58]
  wire  _GEN_423 = 8'ha7 == _T_1[7:0] ? content_167 : _GEN_422; // @[Cat.scala 29:58]
  wire  _GEN_424 = 8'ha8 == _T_1[7:0] ? content_168 : _GEN_423; // @[Cat.scala 29:58]
  wire  _GEN_425 = 8'ha9 == _T_1[7:0] ? content_169 : _GEN_424; // @[Cat.scala 29:58]
  wire  _GEN_426 = 8'haa == _T_1[7:0] ? content_170 : _GEN_425; // @[Cat.scala 29:58]
  wire  _GEN_427 = 8'hab == _T_1[7:0] ? content_171 : _GEN_426; // @[Cat.scala 29:58]
  wire  _GEN_428 = 8'hac == _T_1[7:0] ? content_172 : _GEN_427; // @[Cat.scala 29:58]
  wire  _GEN_429 = 8'had == _T_1[7:0] ? content_173 : _GEN_428; // @[Cat.scala 29:58]
  wire  _GEN_430 = 8'hae == _T_1[7:0] ? content_174 : _GEN_429; // @[Cat.scala 29:58]
  wire  _GEN_431 = 8'haf == _T_1[7:0] ? content_175 : _GEN_430; // @[Cat.scala 29:58]
  wire  _GEN_432 = 8'hb0 == _T_1[7:0] ? content_176 : _GEN_431; // @[Cat.scala 29:58]
  wire  _GEN_433 = 8'hb1 == _T_1[7:0] ? content_177 : _GEN_432; // @[Cat.scala 29:58]
  wire  _GEN_434 = 8'hb2 == _T_1[7:0] ? content_178 : _GEN_433; // @[Cat.scala 29:58]
  wire  _GEN_435 = 8'hb3 == _T_1[7:0] ? content_179 : _GEN_434; // @[Cat.scala 29:58]
  wire  _GEN_436 = 8'hb4 == _T_1[7:0] ? content_180 : _GEN_435; // @[Cat.scala 29:58]
  wire  _GEN_437 = 8'hb5 == _T_1[7:0] ? content_181 : _GEN_436; // @[Cat.scala 29:58]
  wire  _GEN_438 = 8'hb6 == _T_1[7:0] ? content_182 : _GEN_437; // @[Cat.scala 29:58]
  wire  _GEN_439 = 8'hb7 == _T_1[7:0] ? content_183 : _GEN_438; // @[Cat.scala 29:58]
  wire  _GEN_440 = 8'hb8 == _T_1[7:0] ? content_184 : _GEN_439; // @[Cat.scala 29:58]
  wire  _GEN_441 = 8'hb9 == _T_1[7:0] ? content_185 : _GEN_440; // @[Cat.scala 29:58]
  wire  _GEN_442 = 8'hba == _T_1[7:0] ? content_186 : _GEN_441; // @[Cat.scala 29:58]
  wire  _GEN_443 = 8'hbb == _T_1[7:0] ? content_187 : _GEN_442; // @[Cat.scala 29:58]
  wire  _GEN_444 = 8'hbc == _T_1[7:0] ? content_188 : _GEN_443; // @[Cat.scala 29:58]
  wire  _GEN_445 = 8'hbd == _T_1[7:0] ? content_189 : _GEN_444; // @[Cat.scala 29:58]
  wire  _GEN_446 = 8'hbe == _T_1[7:0] ? content_190 : _GEN_445; // @[Cat.scala 29:58]
  wire  _GEN_447 = 8'hbf == _T_1[7:0] ? content_191 : _GEN_446; // @[Cat.scala 29:58]
  wire  _GEN_448 = 8'hc0 == _T_1[7:0] ? content_192 : _GEN_447; // @[Cat.scala 29:58]
  wire  _GEN_449 = 8'hc1 == _T_1[7:0] ? content_193 : _GEN_448; // @[Cat.scala 29:58]
  wire  _GEN_450 = 8'hc2 == _T_1[7:0] ? content_194 : _GEN_449; // @[Cat.scala 29:58]
  wire  _GEN_451 = 8'hc3 == _T_1[7:0] ? content_195 : _GEN_450; // @[Cat.scala 29:58]
  wire  _GEN_452 = 8'hc4 == _T_1[7:0] ? content_196 : _GEN_451; // @[Cat.scala 29:58]
  wire  _GEN_453 = 8'hc5 == _T_1[7:0] ? content_197 : _GEN_452; // @[Cat.scala 29:58]
  wire  _GEN_454 = 8'hc6 == _T_1[7:0] ? content_198 : _GEN_453; // @[Cat.scala 29:58]
  wire  _GEN_455 = 8'hc7 == _T_1[7:0] ? content_199 : _GEN_454; // @[Cat.scala 29:58]
  wire  _GEN_456 = 8'hc8 == _T_1[7:0] ? content_200 : _GEN_455; // @[Cat.scala 29:58]
  wire  _GEN_457 = 8'hc9 == _T_1[7:0] ? content_201 : _GEN_456; // @[Cat.scala 29:58]
  wire  _GEN_458 = 8'hca == _T_1[7:0] ? content_202 : _GEN_457; // @[Cat.scala 29:58]
  wire  _GEN_459 = 8'hcb == _T_1[7:0] ? content_203 : _GEN_458; // @[Cat.scala 29:58]
  wire  _GEN_460 = 8'hcc == _T_1[7:0] ? content_204 : _GEN_459; // @[Cat.scala 29:58]
  wire  _GEN_461 = 8'hcd == _T_1[7:0] ? content_205 : _GEN_460; // @[Cat.scala 29:58]
  wire  _GEN_462 = 8'hce == _T_1[7:0] ? content_206 : _GEN_461; // @[Cat.scala 29:58]
  wire  _GEN_463 = 8'hcf == _T_1[7:0] ? content_207 : _GEN_462; // @[Cat.scala 29:58]
  wire  _GEN_464 = 8'hd0 == _T_1[7:0] ? content_208 : _GEN_463; // @[Cat.scala 29:58]
  wire  _GEN_465 = 8'hd1 == _T_1[7:0] ? content_209 : _GEN_464; // @[Cat.scala 29:58]
  wire  _GEN_466 = 8'hd2 == _T_1[7:0] ? content_210 : _GEN_465; // @[Cat.scala 29:58]
  wire  _GEN_467 = 8'hd3 == _T_1[7:0] ? content_211 : _GEN_466; // @[Cat.scala 29:58]
  wire  _GEN_468 = 8'hd4 == _T_1[7:0] ? content_212 : _GEN_467; // @[Cat.scala 29:58]
  wire  _GEN_469 = 8'hd5 == _T_1[7:0] ? content_213 : _GEN_468; // @[Cat.scala 29:58]
  wire  _GEN_470 = 8'hd6 == _T_1[7:0] ? content_214 : _GEN_469; // @[Cat.scala 29:58]
  wire  _GEN_471 = 8'hd7 == _T_1[7:0] ? content_215 : _GEN_470; // @[Cat.scala 29:58]
  wire  _GEN_472 = 8'hd8 == _T_1[7:0] ? content_216 : _GEN_471; // @[Cat.scala 29:58]
  wire  _GEN_473 = 8'hd9 == _T_1[7:0] ? content_217 : _GEN_472; // @[Cat.scala 29:58]
  wire  _GEN_474 = 8'hda == _T_1[7:0] ? content_218 : _GEN_473; // @[Cat.scala 29:58]
  wire  _GEN_475 = 8'hdb == _T_1[7:0] ? content_219 : _GEN_474; // @[Cat.scala 29:58]
  wire  _GEN_476 = 8'hdc == _T_1[7:0] ? content_220 : _GEN_475; // @[Cat.scala 29:58]
  wire  _GEN_477 = 8'hdd == _T_1[7:0] ? content_221 : _GEN_476; // @[Cat.scala 29:58]
  wire  _GEN_478 = 8'hde == _T_1[7:0] ? content_222 : _GEN_477; // @[Cat.scala 29:58]
  wire  _GEN_479 = 8'hdf == _T_1[7:0] ? content_223 : _GEN_478; // @[Cat.scala 29:58]
  wire  _GEN_480 = 8'he0 == _T_1[7:0] ? content_224 : _GEN_479; // @[Cat.scala 29:58]
  wire  _GEN_481 = 8'he1 == _T_1[7:0] ? content_225 : _GEN_480; // @[Cat.scala 29:58]
  wire  _GEN_482 = 8'he2 == _T_1[7:0] ? content_226 : _GEN_481; // @[Cat.scala 29:58]
  wire  _GEN_483 = 8'he3 == _T_1[7:0] ? content_227 : _GEN_482; // @[Cat.scala 29:58]
  wire  _GEN_484 = 8'he4 == _T_1[7:0] ? content_228 : _GEN_483; // @[Cat.scala 29:58]
  wire  _GEN_485 = 8'he5 == _T_1[7:0] ? content_229 : _GEN_484; // @[Cat.scala 29:58]
  wire  _GEN_486 = 8'he6 == _T_1[7:0] ? content_230 : _GEN_485; // @[Cat.scala 29:58]
  wire  _GEN_487 = 8'he7 == _T_1[7:0] ? content_231 : _GEN_486; // @[Cat.scala 29:58]
  wire  _GEN_488 = 8'he8 == _T_1[7:0] ? content_232 : _GEN_487; // @[Cat.scala 29:58]
  wire  _GEN_489 = 8'he9 == _T_1[7:0] ? content_233 : _GEN_488; // @[Cat.scala 29:58]
  wire  _GEN_490 = 8'hea == _T_1[7:0] ? content_234 : _GEN_489; // @[Cat.scala 29:58]
  wire  _GEN_491 = 8'heb == _T_1[7:0] ? content_235 : _GEN_490; // @[Cat.scala 29:58]
  wire  _GEN_492 = 8'hec == _T_1[7:0] ? content_236 : _GEN_491; // @[Cat.scala 29:58]
  wire  _GEN_493 = 8'hed == _T_1[7:0] ? content_237 : _GEN_492; // @[Cat.scala 29:58]
  wire  _GEN_494 = 8'hee == _T_1[7:0] ? content_238 : _GEN_493; // @[Cat.scala 29:58]
  wire  _GEN_495 = 8'hef == _T_1[7:0] ? content_239 : _GEN_494; // @[Cat.scala 29:58]
  wire  _GEN_496 = 8'hf0 == _T_1[7:0] ? content_240 : _GEN_495; // @[Cat.scala 29:58]
  wire  _GEN_497 = 8'hf1 == _T_1[7:0] ? content_241 : _GEN_496; // @[Cat.scala 29:58]
  wire  _GEN_498 = 8'hf2 == _T_1[7:0] ? content_242 : _GEN_497; // @[Cat.scala 29:58]
  wire  _GEN_499 = 8'hf3 == _T_1[7:0] ? content_243 : _GEN_498; // @[Cat.scala 29:58]
  wire  _GEN_500 = 8'hf4 == _T_1[7:0] ? content_244 : _GEN_499; // @[Cat.scala 29:58]
  wire  _GEN_501 = 8'hf5 == _T_1[7:0] ? content_245 : _GEN_500; // @[Cat.scala 29:58]
  wire  _GEN_502 = 8'hf6 == _T_1[7:0] ? content_246 : _GEN_501; // @[Cat.scala 29:58]
  wire  _GEN_503 = 8'hf7 == _T_1[7:0] ? content_247 : _GEN_502; // @[Cat.scala 29:58]
  wire  _GEN_504 = 8'hf8 == _T_1[7:0] ? content_248 : _GEN_503; // @[Cat.scala 29:58]
  wire  _GEN_505 = 8'hf9 == _T_1[7:0] ? content_249 : _GEN_504; // @[Cat.scala 29:58]
  wire  _GEN_506 = 8'hfa == _T_1[7:0] ? content_250 : _GEN_505; // @[Cat.scala 29:58]
  wire  _GEN_507 = 8'hfb == _T_1[7:0] ? content_251 : _GEN_506; // @[Cat.scala 29:58]
  wire  _GEN_508 = 8'hfc == _T_1[7:0] ? content_252 : _GEN_507; // @[Cat.scala 29:58]
  wire  _GEN_509 = 8'hfd == _T_1[7:0] ? content_253 : _GEN_508; // @[Cat.scala 29:58]
  wire  _GEN_510 = 8'hfe == _T_1[7:0] ? content_254 : _GEN_509; // @[Cat.scala 29:58]
  wire  _GEN_511 = 8'hff == _T_1[7:0] ? content_255 : _GEN_510; // @[Cat.scala 29:58]
  wire  _GEN_513 = 8'h1 == _T_11[7:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_514 = 8'h2 == _T_11[7:0] ? content_2 : _GEN_513; // @[Cat.scala 29:58]
  wire  _GEN_515 = 8'h3 == _T_11[7:0] ? content_3 : _GEN_514; // @[Cat.scala 29:58]
  wire  _GEN_516 = 8'h4 == _T_11[7:0] ? content_4 : _GEN_515; // @[Cat.scala 29:58]
  wire  _GEN_517 = 8'h5 == _T_11[7:0] ? content_5 : _GEN_516; // @[Cat.scala 29:58]
  wire  _GEN_518 = 8'h6 == _T_11[7:0] ? content_6 : _GEN_517; // @[Cat.scala 29:58]
  wire  _GEN_519 = 8'h7 == _T_11[7:0] ? content_7 : _GEN_518; // @[Cat.scala 29:58]
  wire  _GEN_520 = 8'h8 == _T_11[7:0] ? content_8 : _GEN_519; // @[Cat.scala 29:58]
  wire  _GEN_521 = 8'h9 == _T_11[7:0] ? content_9 : _GEN_520; // @[Cat.scala 29:58]
  wire  _GEN_522 = 8'ha == _T_11[7:0] ? content_10 : _GEN_521; // @[Cat.scala 29:58]
  wire  _GEN_523 = 8'hb == _T_11[7:0] ? content_11 : _GEN_522; // @[Cat.scala 29:58]
  wire  _GEN_524 = 8'hc == _T_11[7:0] ? content_12 : _GEN_523; // @[Cat.scala 29:58]
  wire  _GEN_525 = 8'hd == _T_11[7:0] ? content_13 : _GEN_524; // @[Cat.scala 29:58]
  wire  _GEN_526 = 8'he == _T_11[7:0] ? content_14 : _GEN_525; // @[Cat.scala 29:58]
  wire  _GEN_527 = 8'hf == _T_11[7:0] ? content_15 : _GEN_526; // @[Cat.scala 29:58]
  wire  _GEN_528 = 8'h10 == _T_11[7:0] ? content_16 : _GEN_527; // @[Cat.scala 29:58]
  wire  _GEN_529 = 8'h11 == _T_11[7:0] ? content_17 : _GEN_528; // @[Cat.scala 29:58]
  wire  _GEN_530 = 8'h12 == _T_11[7:0] ? content_18 : _GEN_529; // @[Cat.scala 29:58]
  wire  _GEN_531 = 8'h13 == _T_11[7:0] ? content_19 : _GEN_530; // @[Cat.scala 29:58]
  wire  _GEN_532 = 8'h14 == _T_11[7:0] ? content_20 : _GEN_531; // @[Cat.scala 29:58]
  wire  _GEN_533 = 8'h15 == _T_11[7:0] ? content_21 : _GEN_532; // @[Cat.scala 29:58]
  wire  _GEN_534 = 8'h16 == _T_11[7:0] ? content_22 : _GEN_533; // @[Cat.scala 29:58]
  wire  _GEN_535 = 8'h17 == _T_11[7:0] ? content_23 : _GEN_534; // @[Cat.scala 29:58]
  wire  _GEN_536 = 8'h18 == _T_11[7:0] ? content_24 : _GEN_535; // @[Cat.scala 29:58]
  wire  _GEN_537 = 8'h19 == _T_11[7:0] ? content_25 : _GEN_536; // @[Cat.scala 29:58]
  wire  _GEN_538 = 8'h1a == _T_11[7:0] ? content_26 : _GEN_537; // @[Cat.scala 29:58]
  wire  _GEN_539 = 8'h1b == _T_11[7:0] ? content_27 : _GEN_538; // @[Cat.scala 29:58]
  wire  _GEN_540 = 8'h1c == _T_11[7:0] ? content_28 : _GEN_539; // @[Cat.scala 29:58]
  wire  _GEN_541 = 8'h1d == _T_11[7:0] ? content_29 : _GEN_540; // @[Cat.scala 29:58]
  wire  _GEN_542 = 8'h1e == _T_11[7:0] ? content_30 : _GEN_541; // @[Cat.scala 29:58]
  wire  _GEN_543 = 8'h1f == _T_11[7:0] ? content_31 : _GEN_542; // @[Cat.scala 29:58]
  wire  _GEN_544 = 8'h20 == _T_11[7:0] ? content_32 : _GEN_543; // @[Cat.scala 29:58]
  wire  _GEN_545 = 8'h21 == _T_11[7:0] ? content_33 : _GEN_544; // @[Cat.scala 29:58]
  wire  _GEN_546 = 8'h22 == _T_11[7:0] ? content_34 : _GEN_545; // @[Cat.scala 29:58]
  wire  _GEN_547 = 8'h23 == _T_11[7:0] ? content_35 : _GEN_546; // @[Cat.scala 29:58]
  wire  _GEN_548 = 8'h24 == _T_11[7:0] ? content_36 : _GEN_547; // @[Cat.scala 29:58]
  wire  _GEN_549 = 8'h25 == _T_11[7:0] ? content_37 : _GEN_548; // @[Cat.scala 29:58]
  wire  _GEN_550 = 8'h26 == _T_11[7:0] ? content_38 : _GEN_549; // @[Cat.scala 29:58]
  wire  _GEN_551 = 8'h27 == _T_11[7:0] ? content_39 : _GEN_550; // @[Cat.scala 29:58]
  wire  _GEN_552 = 8'h28 == _T_11[7:0] ? content_40 : _GEN_551; // @[Cat.scala 29:58]
  wire  _GEN_553 = 8'h29 == _T_11[7:0] ? content_41 : _GEN_552; // @[Cat.scala 29:58]
  wire  _GEN_554 = 8'h2a == _T_11[7:0] ? content_42 : _GEN_553; // @[Cat.scala 29:58]
  wire  _GEN_555 = 8'h2b == _T_11[7:0] ? content_43 : _GEN_554; // @[Cat.scala 29:58]
  wire  _GEN_556 = 8'h2c == _T_11[7:0] ? content_44 : _GEN_555; // @[Cat.scala 29:58]
  wire  _GEN_557 = 8'h2d == _T_11[7:0] ? content_45 : _GEN_556; // @[Cat.scala 29:58]
  wire  _GEN_558 = 8'h2e == _T_11[7:0] ? content_46 : _GEN_557; // @[Cat.scala 29:58]
  wire  _GEN_559 = 8'h2f == _T_11[7:0] ? content_47 : _GEN_558; // @[Cat.scala 29:58]
  wire  _GEN_560 = 8'h30 == _T_11[7:0] ? content_48 : _GEN_559; // @[Cat.scala 29:58]
  wire  _GEN_561 = 8'h31 == _T_11[7:0] ? content_49 : _GEN_560; // @[Cat.scala 29:58]
  wire  _GEN_562 = 8'h32 == _T_11[7:0] ? content_50 : _GEN_561; // @[Cat.scala 29:58]
  wire  _GEN_563 = 8'h33 == _T_11[7:0] ? content_51 : _GEN_562; // @[Cat.scala 29:58]
  wire  _GEN_564 = 8'h34 == _T_11[7:0] ? content_52 : _GEN_563; // @[Cat.scala 29:58]
  wire  _GEN_565 = 8'h35 == _T_11[7:0] ? content_53 : _GEN_564; // @[Cat.scala 29:58]
  wire  _GEN_566 = 8'h36 == _T_11[7:0] ? content_54 : _GEN_565; // @[Cat.scala 29:58]
  wire  _GEN_567 = 8'h37 == _T_11[7:0] ? content_55 : _GEN_566; // @[Cat.scala 29:58]
  wire  _GEN_568 = 8'h38 == _T_11[7:0] ? content_56 : _GEN_567; // @[Cat.scala 29:58]
  wire  _GEN_569 = 8'h39 == _T_11[7:0] ? content_57 : _GEN_568; // @[Cat.scala 29:58]
  wire  _GEN_570 = 8'h3a == _T_11[7:0] ? content_58 : _GEN_569; // @[Cat.scala 29:58]
  wire  _GEN_571 = 8'h3b == _T_11[7:0] ? content_59 : _GEN_570; // @[Cat.scala 29:58]
  wire  _GEN_572 = 8'h3c == _T_11[7:0] ? content_60 : _GEN_571; // @[Cat.scala 29:58]
  wire  _GEN_573 = 8'h3d == _T_11[7:0] ? content_61 : _GEN_572; // @[Cat.scala 29:58]
  wire  _GEN_574 = 8'h3e == _T_11[7:0] ? content_62 : _GEN_573; // @[Cat.scala 29:58]
  wire  _GEN_575 = 8'h3f == _T_11[7:0] ? content_63 : _GEN_574; // @[Cat.scala 29:58]
  wire  _GEN_576 = 8'h40 == _T_11[7:0] ? content_64 : _GEN_575; // @[Cat.scala 29:58]
  wire  _GEN_577 = 8'h41 == _T_11[7:0] ? content_65 : _GEN_576; // @[Cat.scala 29:58]
  wire  _GEN_578 = 8'h42 == _T_11[7:0] ? content_66 : _GEN_577; // @[Cat.scala 29:58]
  wire  _GEN_579 = 8'h43 == _T_11[7:0] ? content_67 : _GEN_578; // @[Cat.scala 29:58]
  wire  _GEN_580 = 8'h44 == _T_11[7:0] ? content_68 : _GEN_579; // @[Cat.scala 29:58]
  wire  _GEN_581 = 8'h45 == _T_11[7:0] ? content_69 : _GEN_580; // @[Cat.scala 29:58]
  wire  _GEN_582 = 8'h46 == _T_11[7:0] ? content_70 : _GEN_581; // @[Cat.scala 29:58]
  wire  _GEN_583 = 8'h47 == _T_11[7:0] ? content_71 : _GEN_582; // @[Cat.scala 29:58]
  wire  _GEN_584 = 8'h48 == _T_11[7:0] ? content_72 : _GEN_583; // @[Cat.scala 29:58]
  wire  _GEN_585 = 8'h49 == _T_11[7:0] ? content_73 : _GEN_584; // @[Cat.scala 29:58]
  wire  _GEN_586 = 8'h4a == _T_11[7:0] ? content_74 : _GEN_585; // @[Cat.scala 29:58]
  wire  _GEN_587 = 8'h4b == _T_11[7:0] ? content_75 : _GEN_586; // @[Cat.scala 29:58]
  wire  _GEN_588 = 8'h4c == _T_11[7:0] ? content_76 : _GEN_587; // @[Cat.scala 29:58]
  wire  _GEN_589 = 8'h4d == _T_11[7:0] ? content_77 : _GEN_588; // @[Cat.scala 29:58]
  wire  _GEN_590 = 8'h4e == _T_11[7:0] ? content_78 : _GEN_589; // @[Cat.scala 29:58]
  wire  _GEN_591 = 8'h4f == _T_11[7:0] ? content_79 : _GEN_590; // @[Cat.scala 29:58]
  wire  _GEN_592 = 8'h50 == _T_11[7:0] ? content_80 : _GEN_591; // @[Cat.scala 29:58]
  wire  _GEN_593 = 8'h51 == _T_11[7:0] ? content_81 : _GEN_592; // @[Cat.scala 29:58]
  wire  _GEN_594 = 8'h52 == _T_11[7:0] ? content_82 : _GEN_593; // @[Cat.scala 29:58]
  wire  _GEN_595 = 8'h53 == _T_11[7:0] ? content_83 : _GEN_594; // @[Cat.scala 29:58]
  wire  _GEN_596 = 8'h54 == _T_11[7:0] ? content_84 : _GEN_595; // @[Cat.scala 29:58]
  wire  _GEN_597 = 8'h55 == _T_11[7:0] ? content_85 : _GEN_596; // @[Cat.scala 29:58]
  wire  _GEN_598 = 8'h56 == _T_11[7:0] ? content_86 : _GEN_597; // @[Cat.scala 29:58]
  wire  _GEN_599 = 8'h57 == _T_11[7:0] ? content_87 : _GEN_598; // @[Cat.scala 29:58]
  wire  _GEN_600 = 8'h58 == _T_11[7:0] ? content_88 : _GEN_599; // @[Cat.scala 29:58]
  wire  _GEN_601 = 8'h59 == _T_11[7:0] ? content_89 : _GEN_600; // @[Cat.scala 29:58]
  wire  _GEN_602 = 8'h5a == _T_11[7:0] ? content_90 : _GEN_601; // @[Cat.scala 29:58]
  wire  _GEN_603 = 8'h5b == _T_11[7:0] ? content_91 : _GEN_602; // @[Cat.scala 29:58]
  wire  _GEN_604 = 8'h5c == _T_11[7:0] ? content_92 : _GEN_603; // @[Cat.scala 29:58]
  wire  _GEN_605 = 8'h5d == _T_11[7:0] ? content_93 : _GEN_604; // @[Cat.scala 29:58]
  wire  _GEN_606 = 8'h5e == _T_11[7:0] ? content_94 : _GEN_605; // @[Cat.scala 29:58]
  wire  _GEN_607 = 8'h5f == _T_11[7:0] ? content_95 : _GEN_606; // @[Cat.scala 29:58]
  wire  _GEN_608 = 8'h60 == _T_11[7:0] ? content_96 : _GEN_607; // @[Cat.scala 29:58]
  wire  _GEN_609 = 8'h61 == _T_11[7:0] ? content_97 : _GEN_608; // @[Cat.scala 29:58]
  wire  _GEN_610 = 8'h62 == _T_11[7:0] ? content_98 : _GEN_609; // @[Cat.scala 29:58]
  wire  _GEN_611 = 8'h63 == _T_11[7:0] ? content_99 : _GEN_610; // @[Cat.scala 29:58]
  wire  _GEN_612 = 8'h64 == _T_11[7:0] ? content_100 : _GEN_611; // @[Cat.scala 29:58]
  wire  _GEN_613 = 8'h65 == _T_11[7:0] ? content_101 : _GEN_612; // @[Cat.scala 29:58]
  wire  _GEN_614 = 8'h66 == _T_11[7:0] ? content_102 : _GEN_613; // @[Cat.scala 29:58]
  wire  _GEN_615 = 8'h67 == _T_11[7:0] ? content_103 : _GEN_614; // @[Cat.scala 29:58]
  wire  _GEN_616 = 8'h68 == _T_11[7:0] ? content_104 : _GEN_615; // @[Cat.scala 29:58]
  wire  _GEN_617 = 8'h69 == _T_11[7:0] ? content_105 : _GEN_616; // @[Cat.scala 29:58]
  wire  _GEN_618 = 8'h6a == _T_11[7:0] ? content_106 : _GEN_617; // @[Cat.scala 29:58]
  wire  _GEN_619 = 8'h6b == _T_11[7:0] ? content_107 : _GEN_618; // @[Cat.scala 29:58]
  wire  _GEN_620 = 8'h6c == _T_11[7:0] ? content_108 : _GEN_619; // @[Cat.scala 29:58]
  wire  _GEN_621 = 8'h6d == _T_11[7:0] ? content_109 : _GEN_620; // @[Cat.scala 29:58]
  wire  _GEN_622 = 8'h6e == _T_11[7:0] ? content_110 : _GEN_621; // @[Cat.scala 29:58]
  wire  _GEN_623 = 8'h6f == _T_11[7:0] ? content_111 : _GEN_622; // @[Cat.scala 29:58]
  wire  _GEN_624 = 8'h70 == _T_11[7:0] ? content_112 : _GEN_623; // @[Cat.scala 29:58]
  wire  _GEN_625 = 8'h71 == _T_11[7:0] ? content_113 : _GEN_624; // @[Cat.scala 29:58]
  wire  _GEN_626 = 8'h72 == _T_11[7:0] ? content_114 : _GEN_625; // @[Cat.scala 29:58]
  wire  _GEN_627 = 8'h73 == _T_11[7:0] ? content_115 : _GEN_626; // @[Cat.scala 29:58]
  wire  _GEN_628 = 8'h74 == _T_11[7:0] ? content_116 : _GEN_627; // @[Cat.scala 29:58]
  wire  _GEN_629 = 8'h75 == _T_11[7:0] ? content_117 : _GEN_628; // @[Cat.scala 29:58]
  wire  _GEN_630 = 8'h76 == _T_11[7:0] ? content_118 : _GEN_629; // @[Cat.scala 29:58]
  wire  _GEN_631 = 8'h77 == _T_11[7:0] ? content_119 : _GEN_630; // @[Cat.scala 29:58]
  wire  _GEN_632 = 8'h78 == _T_11[7:0] ? content_120 : _GEN_631; // @[Cat.scala 29:58]
  wire  _GEN_633 = 8'h79 == _T_11[7:0] ? content_121 : _GEN_632; // @[Cat.scala 29:58]
  wire  _GEN_634 = 8'h7a == _T_11[7:0] ? content_122 : _GEN_633; // @[Cat.scala 29:58]
  wire  _GEN_635 = 8'h7b == _T_11[7:0] ? content_123 : _GEN_634; // @[Cat.scala 29:58]
  wire  _GEN_636 = 8'h7c == _T_11[7:0] ? content_124 : _GEN_635; // @[Cat.scala 29:58]
  wire  _GEN_637 = 8'h7d == _T_11[7:0] ? content_125 : _GEN_636; // @[Cat.scala 29:58]
  wire  _GEN_638 = 8'h7e == _T_11[7:0] ? content_126 : _GEN_637; // @[Cat.scala 29:58]
  wire  _GEN_639 = 8'h7f == _T_11[7:0] ? content_127 : _GEN_638; // @[Cat.scala 29:58]
  wire  _GEN_640 = 8'h80 == _T_11[7:0] ? content_128 : _GEN_639; // @[Cat.scala 29:58]
  wire  _GEN_641 = 8'h81 == _T_11[7:0] ? content_129 : _GEN_640; // @[Cat.scala 29:58]
  wire  _GEN_642 = 8'h82 == _T_11[7:0] ? content_130 : _GEN_641; // @[Cat.scala 29:58]
  wire  _GEN_643 = 8'h83 == _T_11[7:0] ? content_131 : _GEN_642; // @[Cat.scala 29:58]
  wire  _GEN_644 = 8'h84 == _T_11[7:0] ? content_132 : _GEN_643; // @[Cat.scala 29:58]
  wire  _GEN_645 = 8'h85 == _T_11[7:0] ? content_133 : _GEN_644; // @[Cat.scala 29:58]
  wire  _GEN_646 = 8'h86 == _T_11[7:0] ? content_134 : _GEN_645; // @[Cat.scala 29:58]
  wire  _GEN_647 = 8'h87 == _T_11[7:0] ? content_135 : _GEN_646; // @[Cat.scala 29:58]
  wire  _GEN_648 = 8'h88 == _T_11[7:0] ? content_136 : _GEN_647; // @[Cat.scala 29:58]
  wire  _GEN_649 = 8'h89 == _T_11[7:0] ? content_137 : _GEN_648; // @[Cat.scala 29:58]
  wire  _GEN_650 = 8'h8a == _T_11[7:0] ? content_138 : _GEN_649; // @[Cat.scala 29:58]
  wire  _GEN_651 = 8'h8b == _T_11[7:0] ? content_139 : _GEN_650; // @[Cat.scala 29:58]
  wire  _GEN_652 = 8'h8c == _T_11[7:0] ? content_140 : _GEN_651; // @[Cat.scala 29:58]
  wire  _GEN_653 = 8'h8d == _T_11[7:0] ? content_141 : _GEN_652; // @[Cat.scala 29:58]
  wire  _GEN_654 = 8'h8e == _T_11[7:0] ? content_142 : _GEN_653; // @[Cat.scala 29:58]
  wire  _GEN_655 = 8'h8f == _T_11[7:0] ? content_143 : _GEN_654; // @[Cat.scala 29:58]
  wire  _GEN_656 = 8'h90 == _T_11[7:0] ? content_144 : _GEN_655; // @[Cat.scala 29:58]
  wire  _GEN_657 = 8'h91 == _T_11[7:0] ? content_145 : _GEN_656; // @[Cat.scala 29:58]
  wire  _GEN_658 = 8'h92 == _T_11[7:0] ? content_146 : _GEN_657; // @[Cat.scala 29:58]
  wire  _GEN_659 = 8'h93 == _T_11[7:0] ? content_147 : _GEN_658; // @[Cat.scala 29:58]
  wire  _GEN_660 = 8'h94 == _T_11[7:0] ? content_148 : _GEN_659; // @[Cat.scala 29:58]
  wire  _GEN_661 = 8'h95 == _T_11[7:0] ? content_149 : _GEN_660; // @[Cat.scala 29:58]
  wire  _GEN_662 = 8'h96 == _T_11[7:0] ? content_150 : _GEN_661; // @[Cat.scala 29:58]
  wire  _GEN_663 = 8'h97 == _T_11[7:0] ? content_151 : _GEN_662; // @[Cat.scala 29:58]
  wire  _GEN_664 = 8'h98 == _T_11[7:0] ? content_152 : _GEN_663; // @[Cat.scala 29:58]
  wire  _GEN_665 = 8'h99 == _T_11[7:0] ? content_153 : _GEN_664; // @[Cat.scala 29:58]
  wire  _GEN_666 = 8'h9a == _T_11[7:0] ? content_154 : _GEN_665; // @[Cat.scala 29:58]
  wire  _GEN_667 = 8'h9b == _T_11[7:0] ? content_155 : _GEN_666; // @[Cat.scala 29:58]
  wire  _GEN_668 = 8'h9c == _T_11[7:0] ? content_156 : _GEN_667; // @[Cat.scala 29:58]
  wire  _GEN_669 = 8'h9d == _T_11[7:0] ? content_157 : _GEN_668; // @[Cat.scala 29:58]
  wire  _GEN_670 = 8'h9e == _T_11[7:0] ? content_158 : _GEN_669; // @[Cat.scala 29:58]
  wire  _GEN_671 = 8'h9f == _T_11[7:0] ? content_159 : _GEN_670; // @[Cat.scala 29:58]
  wire  _GEN_672 = 8'ha0 == _T_11[7:0] ? content_160 : _GEN_671; // @[Cat.scala 29:58]
  wire  _GEN_673 = 8'ha1 == _T_11[7:0] ? content_161 : _GEN_672; // @[Cat.scala 29:58]
  wire  _GEN_674 = 8'ha2 == _T_11[7:0] ? content_162 : _GEN_673; // @[Cat.scala 29:58]
  wire  _GEN_675 = 8'ha3 == _T_11[7:0] ? content_163 : _GEN_674; // @[Cat.scala 29:58]
  wire  _GEN_676 = 8'ha4 == _T_11[7:0] ? content_164 : _GEN_675; // @[Cat.scala 29:58]
  wire  _GEN_677 = 8'ha5 == _T_11[7:0] ? content_165 : _GEN_676; // @[Cat.scala 29:58]
  wire  _GEN_678 = 8'ha6 == _T_11[7:0] ? content_166 : _GEN_677; // @[Cat.scala 29:58]
  wire  _GEN_679 = 8'ha7 == _T_11[7:0] ? content_167 : _GEN_678; // @[Cat.scala 29:58]
  wire  _GEN_680 = 8'ha8 == _T_11[7:0] ? content_168 : _GEN_679; // @[Cat.scala 29:58]
  wire  _GEN_681 = 8'ha9 == _T_11[7:0] ? content_169 : _GEN_680; // @[Cat.scala 29:58]
  wire  _GEN_682 = 8'haa == _T_11[7:0] ? content_170 : _GEN_681; // @[Cat.scala 29:58]
  wire  _GEN_683 = 8'hab == _T_11[7:0] ? content_171 : _GEN_682; // @[Cat.scala 29:58]
  wire  _GEN_684 = 8'hac == _T_11[7:0] ? content_172 : _GEN_683; // @[Cat.scala 29:58]
  wire  _GEN_685 = 8'had == _T_11[7:0] ? content_173 : _GEN_684; // @[Cat.scala 29:58]
  wire  _GEN_686 = 8'hae == _T_11[7:0] ? content_174 : _GEN_685; // @[Cat.scala 29:58]
  wire  _GEN_687 = 8'haf == _T_11[7:0] ? content_175 : _GEN_686; // @[Cat.scala 29:58]
  wire  _GEN_688 = 8'hb0 == _T_11[7:0] ? content_176 : _GEN_687; // @[Cat.scala 29:58]
  wire  _GEN_689 = 8'hb1 == _T_11[7:0] ? content_177 : _GEN_688; // @[Cat.scala 29:58]
  wire  _GEN_690 = 8'hb2 == _T_11[7:0] ? content_178 : _GEN_689; // @[Cat.scala 29:58]
  wire  _GEN_691 = 8'hb3 == _T_11[7:0] ? content_179 : _GEN_690; // @[Cat.scala 29:58]
  wire  _GEN_692 = 8'hb4 == _T_11[7:0] ? content_180 : _GEN_691; // @[Cat.scala 29:58]
  wire  _GEN_693 = 8'hb5 == _T_11[7:0] ? content_181 : _GEN_692; // @[Cat.scala 29:58]
  wire  _GEN_694 = 8'hb6 == _T_11[7:0] ? content_182 : _GEN_693; // @[Cat.scala 29:58]
  wire  _GEN_695 = 8'hb7 == _T_11[7:0] ? content_183 : _GEN_694; // @[Cat.scala 29:58]
  wire  _GEN_696 = 8'hb8 == _T_11[7:0] ? content_184 : _GEN_695; // @[Cat.scala 29:58]
  wire  _GEN_697 = 8'hb9 == _T_11[7:0] ? content_185 : _GEN_696; // @[Cat.scala 29:58]
  wire  _GEN_698 = 8'hba == _T_11[7:0] ? content_186 : _GEN_697; // @[Cat.scala 29:58]
  wire  _GEN_699 = 8'hbb == _T_11[7:0] ? content_187 : _GEN_698; // @[Cat.scala 29:58]
  wire  _GEN_700 = 8'hbc == _T_11[7:0] ? content_188 : _GEN_699; // @[Cat.scala 29:58]
  wire  _GEN_701 = 8'hbd == _T_11[7:0] ? content_189 : _GEN_700; // @[Cat.scala 29:58]
  wire  _GEN_702 = 8'hbe == _T_11[7:0] ? content_190 : _GEN_701; // @[Cat.scala 29:58]
  wire  _GEN_703 = 8'hbf == _T_11[7:0] ? content_191 : _GEN_702; // @[Cat.scala 29:58]
  wire  _GEN_704 = 8'hc0 == _T_11[7:0] ? content_192 : _GEN_703; // @[Cat.scala 29:58]
  wire  _GEN_705 = 8'hc1 == _T_11[7:0] ? content_193 : _GEN_704; // @[Cat.scala 29:58]
  wire  _GEN_706 = 8'hc2 == _T_11[7:0] ? content_194 : _GEN_705; // @[Cat.scala 29:58]
  wire  _GEN_707 = 8'hc3 == _T_11[7:0] ? content_195 : _GEN_706; // @[Cat.scala 29:58]
  wire  _GEN_708 = 8'hc4 == _T_11[7:0] ? content_196 : _GEN_707; // @[Cat.scala 29:58]
  wire  _GEN_709 = 8'hc5 == _T_11[7:0] ? content_197 : _GEN_708; // @[Cat.scala 29:58]
  wire  _GEN_710 = 8'hc6 == _T_11[7:0] ? content_198 : _GEN_709; // @[Cat.scala 29:58]
  wire  _GEN_711 = 8'hc7 == _T_11[7:0] ? content_199 : _GEN_710; // @[Cat.scala 29:58]
  wire  _GEN_712 = 8'hc8 == _T_11[7:0] ? content_200 : _GEN_711; // @[Cat.scala 29:58]
  wire  _GEN_713 = 8'hc9 == _T_11[7:0] ? content_201 : _GEN_712; // @[Cat.scala 29:58]
  wire  _GEN_714 = 8'hca == _T_11[7:0] ? content_202 : _GEN_713; // @[Cat.scala 29:58]
  wire  _GEN_715 = 8'hcb == _T_11[7:0] ? content_203 : _GEN_714; // @[Cat.scala 29:58]
  wire  _GEN_716 = 8'hcc == _T_11[7:0] ? content_204 : _GEN_715; // @[Cat.scala 29:58]
  wire  _GEN_717 = 8'hcd == _T_11[7:0] ? content_205 : _GEN_716; // @[Cat.scala 29:58]
  wire  _GEN_718 = 8'hce == _T_11[7:0] ? content_206 : _GEN_717; // @[Cat.scala 29:58]
  wire  _GEN_719 = 8'hcf == _T_11[7:0] ? content_207 : _GEN_718; // @[Cat.scala 29:58]
  wire  _GEN_720 = 8'hd0 == _T_11[7:0] ? content_208 : _GEN_719; // @[Cat.scala 29:58]
  wire  _GEN_721 = 8'hd1 == _T_11[7:0] ? content_209 : _GEN_720; // @[Cat.scala 29:58]
  wire  _GEN_722 = 8'hd2 == _T_11[7:0] ? content_210 : _GEN_721; // @[Cat.scala 29:58]
  wire  _GEN_723 = 8'hd3 == _T_11[7:0] ? content_211 : _GEN_722; // @[Cat.scala 29:58]
  wire  _GEN_724 = 8'hd4 == _T_11[7:0] ? content_212 : _GEN_723; // @[Cat.scala 29:58]
  wire  _GEN_725 = 8'hd5 == _T_11[7:0] ? content_213 : _GEN_724; // @[Cat.scala 29:58]
  wire  _GEN_726 = 8'hd6 == _T_11[7:0] ? content_214 : _GEN_725; // @[Cat.scala 29:58]
  wire  _GEN_727 = 8'hd7 == _T_11[7:0] ? content_215 : _GEN_726; // @[Cat.scala 29:58]
  wire  _GEN_728 = 8'hd8 == _T_11[7:0] ? content_216 : _GEN_727; // @[Cat.scala 29:58]
  wire  _GEN_729 = 8'hd9 == _T_11[7:0] ? content_217 : _GEN_728; // @[Cat.scala 29:58]
  wire  _GEN_730 = 8'hda == _T_11[7:0] ? content_218 : _GEN_729; // @[Cat.scala 29:58]
  wire  _GEN_731 = 8'hdb == _T_11[7:0] ? content_219 : _GEN_730; // @[Cat.scala 29:58]
  wire  _GEN_732 = 8'hdc == _T_11[7:0] ? content_220 : _GEN_731; // @[Cat.scala 29:58]
  wire  _GEN_733 = 8'hdd == _T_11[7:0] ? content_221 : _GEN_732; // @[Cat.scala 29:58]
  wire  _GEN_734 = 8'hde == _T_11[7:0] ? content_222 : _GEN_733; // @[Cat.scala 29:58]
  wire  _GEN_735 = 8'hdf == _T_11[7:0] ? content_223 : _GEN_734; // @[Cat.scala 29:58]
  wire  _GEN_736 = 8'he0 == _T_11[7:0] ? content_224 : _GEN_735; // @[Cat.scala 29:58]
  wire  _GEN_737 = 8'he1 == _T_11[7:0] ? content_225 : _GEN_736; // @[Cat.scala 29:58]
  wire  _GEN_738 = 8'he2 == _T_11[7:0] ? content_226 : _GEN_737; // @[Cat.scala 29:58]
  wire  _GEN_739 = 8'he3 == _T_11[7:0] ? content_227 : _GEN_738; // @[Cat.scala 29:58]
  wire  _GEN_740 = 8'he4 == _T_11[7:0] ? content_228 : _GEN_739; // @[Cat.scala 29:58]
  wire  _GEN_741 = 8'he5 == _T_11[7:0] ? content_229 : _GEN_740; // @[Cat.scala 29:58]
  wire  _GEN_742 = 8'he6 == _T_11[7:0] ? content_230 : _GEN_741; // @[Cat.scala 29:58]
  wire  _GEN_743 = 8'he7 == _T_11[7:0] ? content_231 : _GEN_742; // @[Cat.scala 29:58]
  wire  _GEN_744 = 8'he8 == _T_11[7:0] ? content_232 : _GEN_743; // @[Cat.scala 29:58]
  wire  _GEN_745 = 8'he9 == _T_11[7:0] ? content_233 : _GEN_744; // @[Cat.scala 29:58]
  wire  _GEN_746 = 8'hea == _T_11[7:0] ? content_234 : _GEN_745; // @[Cat.scala 29:58]
  wire  _GEN_747 = 8'heb == _T_11[7:0] ? content_235 : _GEN_746; // @[Cat.scala 29:58]
  wire  _GEN_748 = 8'hec == _T_11[7:0] ? content_236 : _GEN_747; // @[Cat.scala 29:58]
  wire  _GEN_749 = 8'hed == _T_11[7:0] ? content_237 : _GEN_748; // @[Cat.scala 29:58]
  wire  _GEN_750 = 8'hee == _T_11[7:0] ? content_238 : _GEN_749; // @[Cat.scala 29:58]
  wire  _GEN_751 = 8'hef == _T_11[7:0] ? content_239 : _GEN_750; // @[Cat.scala 29:58]
  wire  _GEN_752 = 8'hf0 == _T_11[7:0] ? content_240 : _GEN_751; // @[Cat.scala 29:58]
  wire  _GEN_753 = 8'hf1 == _T_11[7:0] ? content_241 : _GEN_752; // @[Cat.scala 29:58]
  wire  _GEN_754 = 8'hf2 == _T_11[7:0] ? content_242 : _GEN_753; // @[Cat.scala 29:58]
  wire  _GEN_755 = 8'hf3 == _T_11[7:0] ? content_243 : _GEN_754; // @[Cat.scala 29:58]
  wire  _GEN_756 = 8'hf4 == _T_11[7:0] ? content_244 : _GEN_755; // @[Cat.scala 29:58]
  wire  _GEN_757 = 8'hf5 == _T_11[7:0] ? content_245 : _GEN_756; // @[Cat.scala 29:58]
  wire  _GEN_758 = 8'hf6 == _T_11[7:0] ? content_246 : _GEN_757; // @[Cat.scala 29:58]
  wire  _GEN_759 = 8'hf7 == _T_11[7:0] ? content_247 : _GEN_758; // @[Cat.scala 29:58]
  wire  _GEN_760 = 8'hf8 == _T_11[7:0] ? content_248 : _GEN_759; // @[Cat.scala 29:58]
  wire  _GEN_761 = 8'hf9 == _T_11[7:0] ? content_249 : _GEN_760; // @[Cat.scala 29:58]
  wire  _GEN_762 = 8'hfa == _T_11[7:0] ? content_250 : _GEN_761; // @[Cat.scala 29:58]
  wire  _GEN_763 = 8'hfb == _T_11[7:0] ? content_251 : _GEN_762; // @[Cat.scala 29:58]
  wire  _GEN_764 = 8'hfc == _T_11[7:0] ? content_252 : _GEN_763; // @[Cat.scala 29:58]
  wire  _GEN_765 = 8'hfd == _T_11[7:0] ? content_253 : _GEN_764; // @[Cat.scala 29:58]
  wire  _GEN_766 = 8'hfe == _T_11[7:0] ? content_254 : _GEN_765; // @[Cat.scala 29:58]
  wire  _GEN_767 = 8'hff == _T_11[7:0] ? content_255 : _GEN_766; // @[Cat.scala 29:58]
  wire  _GEN_769 = 8'h1 == _T_8[7:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_770 = 8'h2 == _T_8[7:0] ? content_2 : _GEN_769; // @[Cat.scala 29:58]
  wire  _GEN_771 = 8'h3 == _T_8[7:0] ? content_3 : _GEN_770; // @[Cat.scala 29:58]
  wire  _GEN_772 = 8'h4 == _T_8[7:0] ? content_4 : _GEN_771; // @[Cat.scala 29:58]
  wire  _GEN_773 = 8'h5 == _T_8[7:0] ? content_5 : _GEN_772; // @[Cat.scala 29:58]
  wire  _GEN_774 = 8'h6 == _T_8[7:0] ? content_6 : _GEN_773; // @[Cat.scala 29:58]
  wire  _GEN_775 = 8'h7 == _T_8[7:0] ? content_7 : _GEN_774; // @[Cat.scala 29:58]
  wire  _GEN_776 = 8'h8 == _T_8[7:0] ? content_8 : _GEN_775; // @[Cat.scala 29:58]
  wire  _GEN_777 = 8'h9 == _T_8[7:0] ? content_9 : _GEN_776; // @[Cat.scala 29:58]
  wire  _GEN_778 = 8'ha == _T_8[7:0] ? content_10 : _GEN_777; // @[Cat.scala 29:58]
  wire  _GEN_779 = 8'hb == _T_8[7:0] ? content_11 : _GEN_778; // @[Cat.scala 29:58]
  wire  _GEN_780 = 8'hc == _T_8[7:0] ? content_12 : _GEN_779; // @[Cat.scala 29:58]
  wire  _GEN_781 = 8'hd == _T_8[7:0] ? content_13 : _GEN_780; // @[Cat.scala 29:58]
  wire  _GEN_782 = 8'he == _T_8[7:0] ? content_14 : _GEN_781; // @[Cat.scala 29:58]
  wire  _GEN_783 = 8'hf == _T_8[7:0] ? content_15 : _GEN_782; // @[Cat.scala 29:58]
  wire  _GEN_784 = 8'h10 == _T_8[7:0] ? content_16 : _GEN_783; // @[Cat.scala 29:58]
  wire  _GEN_785 = 8'h11 == _T_8[7:0] ? content_17 : _GEN_784; // @[Cat.scala 29:58]
  wire  _GEN_786 = 8'h12 == _T_8[7:0] ? content_18 : _GEN_785; // @[Cat.scala 29:58]
  wire  _GEN_787 = 8'h13 == _T_8[7:0] ? content_19 : _GEN_786; // @[Cat.scala 29:58]
  wire  _GEN_788 = 8'h14 == _T_8[7:0] ? content_20 : _GEN_787; // @[Cat.scala 29:58]
  wire  _GEN_789 = 8'h15 == _T_8[7:0] ? content_21 : _GEN_788; // @[Cat.scala 29:58]
  wire  _GEN_790 = 8'h16 == _T_8[7:0] ? content_22 : _GEN_789; // @[Cat.scala 29:58]
  wire  _GEN_791 = 8'h17 == _T_8[7:0] ? content_23 : _GEN_790; // @[Cat.scala 29:58]
  wire  _GEN_792 = 8'h18 == _T_8[7:0] ? content_24 : _GEN_791; // @[Cat.scala 29:58]
  wire  _GEN_793 = 8'h19 == _T_8[7:0] ? content_25 : _GEN_792; // @[Cat.scala 29:58]
  wire  _GEN_794 = 8'h1a == _T_8[7:0] ? content_26 : _GEN_793; // @[Cat.scala 29:58]
  wire  _GEN_795 = 8'h1b == _T_8[7:0] ? content_27 : _GEN_794; // @[Cat.scala 29:58]
  wire  _GEN_796 = 8'h1c == _T_8[7:0] ? content_28 : _GEN_795; // @[Cat.scala 29:58]
  wire  _GEN_797 = 8'h1d == _T_8[7:0] ? content_29 : _GEN_796; // @[Cat.scala 29:58]
  wire  _GEN_798 = 8'h1e == _T_8[7:0] ? content_30 : _GEN_797; // @[Cat.scala 29:58]
  wire  _GEN_799 = 8'h1f == _T_8[7:0] ? content_31 : _GEN_798; // @[Cat.scala 29:58]
  wire  _GEN_800 = 8'h20 == _T_8[7:0] ? content_32 : _GEN_799; // @[Cat.scala 29:58]
  wire  _GEN_801 = 8'h21 == _T_8[7:0] ? content_33 : _GEN_800; // @[Cat.scala 29:58]
  wire  _GEN_802 = 8'h22 == _T_8[7:0] ? content_34 : _GEN_801; // @[Cat.scala 29:58]
  wire  _GEN_803 = 8'h23 == _T_8[7:0] ? content_35 : _GEN_802; // @[Cat.scala 29:58]
  wire  _GEN_804 = 8'h24 == _T_8[7:0] ? content_36 : _GEN_803; // @[Cat.scala 29:58]
  wire  _GEN_805 = 8'h25 == _T_8[7:0] ? content_37 : _GEN_804; // @[Cat.scala 29:58]
  wire  _GEN_806 = 8'h26 == _T_8[7:0] ? content_38 : _GEN_805; // @[Cat.scala 29:58]
  wire  _GEN_807 = 8'h27 == _T_8[7:0] ? content_39 : _GEN_806; // @[Cat.scala 29:58]
  wire  _GEN_808 = 8'h28 == _T_8[7:0] ? content_40 : _GEN_807; // @[Cat.scala 29:58]
  wire  _GEN_809 = 8'h29 == _T_8[7:0] ? content_41 : _GEN_808; // @[Cat.scala 29:58]
  wire  _GEN_810 = 8'h2a == _T_8[7:0] ? content_42 : _GEN_809; // @[Cat.scala 29:58]
  wire  _GEN_811 = 8'h2b == _T_8[7:0] ? content_43 : _GEN_810; // @[Cat.scala 29:58]
  wire  _GEN_812 = 8'h2c == _T_8[7:0] ? content_44 : _GEN_811; // @[Cat.scala 29:58]
  wire  _GEN_813 = 8'h2d == _T_8[7:0] ? content_45 : _GEN_812; // @[Cat.scala 29:58]
  wire  _GEN_814 = 8'h2e == _T_8[7:0] ? content_46 : _GEN_813; // @[Cat.scala 29:58]
  wire  _GEN_815 = 8'h2f == _T_8[7:0] ? content_47 : _GEN_814; // @[Cat.scala 29:58]
  wire  _GEN_816 = 8'h30 == _T_8[7:0] ? content_48 : _GEN_815; // @[Cat.scala 29:58]
  wire  _GEN_817 = 8'h31 == _T_8[7:0] ? content_49 : _GEN_816; // @[Cat.scala 29:58]
  wire  _GEN_818 = 8'h32 == _T_8[7:0] ? content_50 : _GEN_817; // @[Cat.scala 29:58]
  wire  _GEN_819 = 8'h33 == _T_8[7:0] ? content_51 : _GEN_818; // @[Cat.scala 29:58]
  wire  _GEN_820 = 8'h34 == _T_8[7:0] ? content_52 : _GEN_819; // @[Cat.scala 29:58]
  wire  _GEN_821 = 8'h35 == _T_8[7:0] ? content_53 : _GEN_820; // @[Cat.scala 29:58]
  wire  _GEN_822 = 8'h36 == _T_8[7:0] ? content_54 : _GEN_821; // @[Cat.scala 29:58]
  wire  _GEN_823 = 8'h37 == _T_8[7:0] ? content_55 : _GEN_822; // @[Cat.scala 29:58]
  wire  _GEN_824 = 8'h38 == _T_8[7:0] ? content_56 : _GEN_823; // @[Cat.scala 29:58]
  wire  _GEN_825 = 8'h39 == _T_8[7:0] ? content_57 : _GEN_824; // @[Cat.scala 29:58]
  wire  _GEN_826 = 8'h3a == _T_8[7:0] ? content_58 : _GEN_825; // @[Cat.scala 29:58]
  wire  _GEN_827 = 8'h3b == _T_8[7:0] ? content_59 : _GEN_826; // @[Cat.scala 29:58]
  wire  _GEN_828 = 8'h3c == _T_8[7:0] ? content_60 : _GEN_827; // @[Cat.scala 29:58]
  wire  _GEN_829 = 8'h3d == _T_8[7:0] ? content_61 : _GEN_828; // @[Cat.scala 29:58]
  wire  _GEN_830 = 8'h3e == _T_8[7:0] ? content_62 : _GEN_829; // @[Cat.scala 29:58]
  wire  _GEN_831 = 8'h3f == _T_8[7:0] ? content_63 : _GEN_830; // @[Cat.scala 29:58]
  wire  _GEN_832 = 8'h40 == _T_8[7:0] ? content_64 : _GEN_831; // @[Cat.scala 29:58]
  wire  _GEN_833 = 8'h41 == _T_8[7:0] ? content_65 : _GEN_832; // @[Cat.scala 29:58]
  wire  _GEN_834 = 8'h42 == _T_8[7:0] ? content_66 : _GEN_833; // @[Cat.scala 29:58]
  wire  _GEN_835 = 8'h43 == _T_8[7:0] ? content_67 : _GEN_834; // @[Cat.scala 29:58]
  wire  _GEN_836 = 8'h44 == _T_8[7:0] ? content_68 : _GEN_835; // @[Cat.scala 29:58]
  wire  _GEN_837 = 8'h45 == _T_8[7:0] ? content_69 : _GEN_836; // @[Cat.scala 29:58]
  wire  _GEN_838 = 8'h46 == _T_8[7:0] ? content_70 : _GEN_837; // @[Cat.scala 29:58]
  wire  _GEN_839 = 8'h47 == _T_8[7:0] ? content_71 : _GEN_838; // @[Cat.scala 29:58]
  wire  _GEN_840 = 8'h48 == _T_8[7:0] ? content_72 : _GEN_839; // @[Cat.scala 29:58]
  wire  _GEN_841 = 8'h49 == _T_8[7:0] ? content_73 : _GEN_840; // @[Cat.scala 29:58]
  wire  _GEN_842 = 8'h4a == _T_8[7:0] ? content_74 : _GEN_841; // @[Cat.scala 29:58]
  wire  _GEN_843 = 8'h4b == _T_8[7:0] ? content_75 : _GEN_842; // @[Cat.scala 29:58]
  wire  _GEN_844 = 8'h4c == _T_8[7:0] ? content_76 : _GEN_843; // @[Cat.scala 29:58]
  wire  _GEN_845 = 8'h4d == _T_8[7:0] ? content_77 : _GEN_844; // @[Cat.scala 29:58]
  wire  _GEN_846 = 8'h4e == _T_8[7:0] ? content_78 : _GEN_845; // @[Cat.scala 29:58]
  wire  _GEN_847 = 8'h4f == _T_8[7:0] ? content_79 : _GEN_846; // @[Cat.scala 29:58]
  wire  _GEN_848 = 8'h50 == _T_8[7:0] ? content_80 : _GEN_847; // @[Cat.scala 29:58]
  wire  _GEN_849 = 8'h51 == _T_8[7:0] ? content_81 : _GEN_848; // @[Cat.scala 29:58]
  wire  _GEN_850 = 8'h52 == _T_8[7:0] ? content_82 : _GEN_849; // @[Cat.scala 29:58]
  wire  _GEN_851 = 8'h53 == _T_8[7:0] ? content_83 : _GEN_850; // @[Cat.scala 29:58]
  wire  _GEN_852 = 8'h54 == _T_8[7:0] ? content_84 : _GEN_851; // @[Cat.scala 29:58]
  wire  _GEN_853 = 8'h55 == _T_8[7:0] ? content_85 : _GEN_852; // @[Cat.scala 29:58]
  wire  _GEN_854 = 8'h56 == _T_8[7:0] ? content_86 : _GEN_853; // @[Cat.scala 29:58]
  wire  _GEN_855 = 8'h57 == _T_8[7:0] ? content_87 : _GEN_854; // @[Cat.scala 29:58]
  wire  _GEN_856 = 8'h58 == _T_8[7:0] ? content_88 : _GEN_855; // @[Cat.scala 29:58]
  wire  _GEN_857 = 8'h59 == _T_8[7:0] ? content_89 : _GEN_856; // @[Cat.scala 29:58]
  wire  _GEN_858 = 8'h5a == _T_8[7:0] ? content_90 : _GEN_857; // @[Cat.scala 29:58]
  wire  _GEN_859 = 8'h5b == _T_8[7:0] ? content_91 : _GEN_858; // @[Cat.scala 29:58]
  wire  _GEN_860 = 8'h5c == _T_8[7:0] ? content_92 : _GEN_859; // @[Cat.scala 29:58]
  wire  _GEN_861 = 8'h5d == _T_8[7:0] ? content_93 : _GEN_860; // @[Cat.scala 29:58]
  wire  _GEN_862 = 8'h5e == _T_8[7:0] ? content_94 : _GEN_861; // @[Cat.scala 29:58]
  wire  _GEN_863 = 8'h5f == _T_8[7:0] ? content_95 : _GEN_862; // @[Cat.scala 29:58]
  wire  _GEN_864 = 8'h60 == _T_8[7:0] ? content_96 : _GEN_863; // @[Cat.scala 29:58]
  wire  _GEN_865 = 8'h61 == _T_8[7:0] ? content_97 : _GEN_864; // @[Cat.scala 29:58]
  wire  _GEN_866 = 8'h62 == _T_8[7:0] ? content_98 : _GEN_865; // @[Cat.scala 29:58]
  wire  _GEN_867 = 8'h63 == _T_8[7:0] ? content_99 : _GEN_866; // @[Cat.scala 29:58]
  wire  _GEN_868 = 8'h64 == _T_8[7:0] ? content_100 : _GEN_867; // @[Cat.scala 29:58]
  wire  _GEN_869 = 8'h65 == _T_8[7:0] ? content_101 : _GEN_868; // @[Cat.scala 29:58]
  wire  _GEN_870 = 8'h66 == _T_8[7:0] ? content_102 : _GEN_869; // @[Cat.scala 29:58]
  wire  _GEN_871 = 8'h67 == _T_8[7:0] ? content_103 : _GEN_870; // @[Cat.scala 29:58]
  wire  _GEN_872 = 8'h68 == _T_8[7:0] ? content_104 : _GEN_871; // @[Cat.scala 29:58]
  wire  _GEN_873 = 8'h69 == _T_8[7:0] ? content_105 : _GEN_872; // @[Cat.scala 29:58]
  wire  _GEN_874 = 8'h6a == _T_8[7:0] ? content_106 : _GEN_873; // @[Cat.scala 29:58]
  wire  _GEN_875 = 8'h6b == _T_8[7:0] ? content_107 : _GEN_874; // @[Cat.scala 29:58]
  wire  _GEN_876 = 8'h6c == _T_8[7:0] ? content_108 : _GEN_875; // @[Cat.scala 29:58]
  wire  _GEN_877 = 8'h6d == _T_8[7:0] ? content_109 : _GEN_876; // @[Cat.scala 29:58]
  wire  _GEN_878 = 8'h6e == _T_8[7:0] ? content_110 : _GEN_877; // @[Cat.scala 29:58]
  wire  _GEN_879 = 8'h6f == _T_8[7:0] ? content_111 : _GEN_878; // @[Cat.scala 29:58]
  wire  _GEN_880 = 8'h70 == _T_8[7:0] ? content_112 : _GEN_879; // @[Cat.scala 29:58]
  wire  _GEN_881 = 8'h71 == _T_8[7:0] ? content_113 : _GEN_880; // @[Cat.scala 29:58]
  wire  _GEN_882 = 8'h72 == _T_8[7:0] ? content_114 : _GEN_881; // @[Cat.scala 29:58]
  wire  _GEN_883 = 8'h73 == _T_8[7:0] ? content_115 : _GEN_882; // @[Cat.scala 29:58]
  wire  _GEN_884 = 8'h74 == _T_8[7:0] ? content_116 : _GEN_883; // @[Cat.scala 29:58]
  wire  _GEN_885 = 8'h75 == _T_8[7:0] ? content_117 : _GEN_884; // @[Cat.scala 29:58]
  wire  _GEN_886 = 8'h76 == _T_8[7:0] ? content_118 : _GEN_885; // @[Cat.scala 29:58]
  wire  _GEN_887 = 8'h77 == _T_8[7:0] ? content_119 : _GEN_886; // @[Cat.scala 29:58]
  wire  _GEN_888 = 8'h78 == _T_8[7:0] ? content_120 : _GEN_887; // @[Cat.scala 29:58]
  wire  _GEN_889 = 8'h79 == _T_8[7:0] ? content_121 : _GEN_888; // @[Cat.scala 29:58]
  wire  _GEN_890 = 8'h7a == _T_8[7:0] ? content_122 : _GEN_889; // @[Cat.scala 29:58]
  wire  _GEN_891 = 8'h7b == _T_8[7:0] ? content_123 : _GEN_890; // @[Cat.scala 29:58]
  wire  _GEN_892 = 8'h7c == _T_8[7:0] ? content_124 : _GEN_891; // @[Cat.scala 29:58]
  wire  _GEN_893 = 8'h7d == _T_8[7:0] ? content_125 : _GEN_892; // @[Cat.scala 29:58]
  wire  _GEN_894 = 8'h7e == _T_8[7:0] ? content_126 : _GEN_893; // @[Cat.scala 29:58]
  wire  _GEN_895 = 8'h7f == _T_8[7:0] ? content_127 : _GEN_894; // @[Cat.scala 29:58]
  wire  _GEN_896 = 8'h80 == _T_8[7:0] ? content_128 : _GEN_895; // @[Cat.scala 29:58]
  wire  _GEN_897 = 8'h81 == _T_8[7:0] ? content_129 : _GEN_896; // @[Cat.scala 29:58]
  wire  _GEN_898 = 8'h82 == _T_8[7:0] ? content_130 : _GEN_897; // @[Cat.scala 29:58]
  wire  _GEN_899 = 8'h83 == _T_8[7:0] ? content_131 : _GEN_898; // @[Cat.scala 29:58]
  wire  _GEN_900 = 8'h84 == _T_8[7:0] ? content_132 : _GEN_899; // @[Cat.scala 29:58]
  wire  _GEN_901 = 8'h85 == _T_8[7:0] ? content_133 : _GEN_900; // @[Cat.scala 29:58]
  wire  _GEN_902 = 8'h86 == _T_8[7:0] ? content_134 : _GEN_901; // @[Cat.scala 29:58]
  wire  _GEN_903 = 8'h87 == _T_8[7:0] ? content_135 : _GEN_902; // @[Cat.scala 29:58]
  wire  _GEN_904 = 8'h88 == _T_8[7:0] ? content_136 : _GEN_903; // @[Cat.scala 29:58]
  wire  _GEN_905 = 8'h89 == _T_8[7:0] ? content_137 : _GEN_904; // @[Cat.scala 29:58]
  wire  _GEN_906 = 8'h8a == _T_8[7:0] ? content_138 : _GEN_905; // @[Cat.scala 29:58]
  wire  _GEN_907 = 8'h8b == _T_8[7:0] ? content_139 : _GEN_906; // @[Cat.scala 29:58]
  wire  _GEN_908 = 8'h8c == _T_8[7:0] ? content_140 : _GEN_907; // @[Cat.scala 29:58]
  wire  _GEN_909 = 8'h8d == _T_8[7:0] ? content_141 : _GEN_908; // @[Cat.scala 29:58]
  wire  _GEN_910 = 8'h8e == _T_8[7:0] ? content_142 : _GEN_909; // @[Cat.scala 29:58]
  wire  _GEN_911 = 8'h8f == _T_8[7:0] ? content_143 : _GEN_910; // @[Cat.scala 29:58]
  wire  _GEN_912 = 8'h90 == _T_8[7:0] ? content_144 : _GEN_911; // @[Cat.scala 29:58]
  wire  _GEN_913 = 8'h91 == _T_8[7:0] ? content_145 : _GEN_912; // @[Cat.scala 29:58]
  wire  _GEN_914 = 8'h92 == _T_8[7:0] ? content_146 : _GEN_913; // @[Cat.scala 29:58]
  wire  _GEN_915 = 8'h93 == _T_8[7:0] ? content_147 : _GEN_914; // @[Cat.scala 29:58]
  wire  _GEN_916 = 8'h94 == _T_8[7:0] ? content_148 : _GEN_915; // @[Cat.scala 29:58]
  wire  _GEN_917 = 8'h95 == _T_8[7:0] ? content_149 : _GEN_916; // @[Cat.scala 29:58]
  wire  _GEN_918 = 8'h96 == _T_8[7:0] ? content_150 : _GEN_917; // @[Cat.scala 29:58]
  wire  _GEN_919 = 8'h97 == _T_8[7:0] ? content_151 : _GEN_918; // @[Cat.scala 29:58]
  wire  _GEN_920 = 8'h98 == _T_8[7:0] ? content_152 : _GEN_919; // @[Cat.scala 29:58]
  wire  _GEN_921 = 8'h99 == _T_8[7:0] ? content_153 : _GEN_920; // @[Cat.scala 29:58]
  wire  _GEN_922 = 8'h9a == _T_8[7:0] ? content_154 : _GEN_921; // @[Cat.scala 29:58]
  wire  _GEN_923 = 8'h9b == _T_8[7:0] ? content_155 : _GEN_922; // @[Cat.scala 29:58]
  wire  _GEN_924 = 8'h9c == _T_8[7:0] ? content_156 : _GEN_923; // @[Cat.scala 29:58]
  wire  _GEN_925 = 8'h9d == _T_8[7:0] ? content_157 : _GEN_924; // @[Cat.scala 29:58]
  wire  _GEN_926 = 8'h9e == _T_8[7:0] ? content_158 : _GEN_925; // @[Cat.scala 29:58]
  wire  _GEN_927 = 8'h9f == _T_8[7:0] ? content_159 : _GEN_926; // @[Cat.scala 29:58]
  wire  _GEN_928 = 8'ha0 == _T_8[7:0] ? content_160 : _GEN_927; // @[Cat.scala 29:58]
  wire  _GEN_929 = 8'ha1 == _T_8[7:0] ? content_161 : _GEN_928; // @[Cat.scala 29:58]
  wire  _GEN_930 = 8'ha2 == _T_8[7:0] ? content_162 : _GEN_929; // @[Cat.scala 29:58]
  wire  _GEN_931 = 8'ha3 == _T_8[7:0] ? content_163 : _GEN_930; // @[Cat.scala 29:58]
  wire  _GEN_932 = 8'ha4 == _T_8[7:0] ? content_164 : _GEN_931; // @[Cat.scala 29:58]
  wire  _GEN_933 = 8'ha5 == _T_8[7:0] ? content_165 : _GEN_932; // @[Cat.scala 29:58]
  wire  _GEN_934 = 8'ha6 == _T_8[7:0] ? content_166 : _GEN_933; // @[Cat.scala 29:58]
  wire  _GEN_935 = 8'ha7 == _T_8[7:0] ? content_167 : _GEN_934; // @[Cat.scala 29:58]
  wire  _GEN_936 = 8'ha8 == _T_8[7:0] ? content_168 : _GEN_935; // @[Cat.scala 29:58]
  wire  _GEN_937 = 8'ha9 == _T_8[7:0] ? content_169 : _GEN_936; // @[Cat.scala 29:58]
  wire  _GEN_938 = 8'haa == _T_8[7:0] ? content_170 : _GEN_937; // @[Cat.scala 29:58]
  wire  _GEN_939 = 8'hab == _T_8[7:0] ? content_171 : _GEN_938; // @[Cat.scala 29:58]
  wire  _GEN_940 = 8'hac == _T_8[7:0] ? content_172 : _GEN_939; // @[Cat.scala 29:58]
  wire  _GEN_941 = 8'had == _T_8[7:0] ? content_173 : _GEN_940; // @[Cat.scala 29:58]
  wire  _GEN_942 = 8'hae == _T_8[7:0] ? content_174 : _GEN_941; // @[Cat.scala 29:58]
  wire  _GEN_943 = 8'haf == _T_8[7:0] ? content_175 : _GEN_942; // @[Cat.scala 29:58]
  wire  _GEN_944 = 8'hb0 == _T_8[7:0] ? content_176 : _GEN_943; // @[Cat.scala 29:58]
  wire  _GEN_945 = 8'hb1 == _T_8[7:0] ? content_177 : _GEN_944; // @[Cat.scala 29:58]
  wire  _GEN_946 = 8'hb2 == _T_8[7:0] ? content_178 : _GEN_945; // @[Cat.scala 29:58]
  wire  _GEN_947 = 8'hb3 == _T_8[7:0] ? content_179 : _GEN_946; // @[Cat.scala 29:58]
  wire  _GEN_948 = 8'hb4 == _T_8[7:0] ? content_180 : _GEN_947; // @[Cat.scala 29:58]
  wire  _GEN_949 = 8'hb5 == _T_8[7:0] ? content_181 : _GEN_948; // @[Cat.scala 29:58]
  wire  _GEN_950 = 8'hb6 == _T_8[7:0] ? content_182 : _GEN_949; // @[Cat.scala 29:58]
  wire  _GEN_951 = 8'hb7 == _T_8[7:0] ? content_183 : _GEN_950; // @[Cat.scala 29:58]
  wire  _GEN_952 = 8'hb8 == _T_8[7:0] ? content_184 : _GEN_951; // @[Cat.scala 29:58]
  wire  _GEN_953 = 8'hb9 == _T_8[7:0] ? content_185 : _GEN_952; // @[Cat.scala 29:58]
  wire  _GEN_954 = 8'hba == _T_8[7:0] ? content_186 : _GEN_953; // @[Cat.scala 29:58]
  wire  _GEN_955 = 8'hbb == _T_8[7:0] ? content_187 : _GEN_954; // @[Cat.scala 29:58]
  wire  _GEN_956 = 8'hbc == _T_8[7:0] ? content_188 : _GEN_955; // @[Cat.scala 29:58]
  wire  _GEN_957 = 8'hbd == _T_8[7:0] ? content_189 : _GEN_956; // @[Cat.scala 29:58]
  wire  _GEN_958 = 8'hbe == _T_8[7:0] ? content_190 : _GEN_957; // @[Cat.scala 29:58]
  wire  _GEN_959 = 8'hbf == _T_8[7:0] ? content_191 : _GEN_958; // @[Cat.scala 29:58]
  wire  _GEN_960 = 8'hc0 == _T_8[7:0] ? content_192 : _GEN_959; // @[Cat.scala 29:58]
  wire  _GEN_961 = 8'hc1 == _T_8[7:0] ? content_193 : _GEN_960; // @[Cat.scala 29:58]
  wire  _GEN_962 = 8'hc2 == _T_8[7:0] ? content_194 : _GEN_961; // @[Cat.scala 29:58]
  wire  _GEN_963 = 8'hc3 == _T_8[7:0] ? content_195 : _GEN_962; // @[Cat.scala 29:58]
  wire  _GEN_964 = 8'hc4 == _T_8[7:0] ? content_196 : _GEN_963; // @[Cat.scala 29:58]
  wire  _GEN_965 = 8'hc5 == _T_8[7:0] ? content_197 : _GEN_964; // @[Cat.scala 29:58]
  wire  _GEN_966 = 8'hc6 == _T_8[7:0] ? content_198 : _GEN_965; // @[Cat.scala 29:58]
  wire  _GEN_967 = 8'hc7 == _T_8[7:0] ? content_199 : _GEN_966; // @[Cat.scala 29:58]
  wire  _GEN_968 = 8'hc8 == _T_8[7:0] ? content_200 : _GEN_967; // @[Cat.scala 29:58]
  wire  _GEN_969 = 8'hc9 == _T_8[7:0] ? content_201 : _GEN_968; // @[Cat.scala 29:58]
  wire  _GEN_970 = 8'hca == _T_8[7:0] ? content_202 : _GEN_969; // @[Cat.scala 29:58]
  wire  _GEN_971 = 8'hcb == _T_8[7:0] ? content_203 : _GEN_970; // @[Cat.scala 29:58]
  wire  _GEN_972 = 8'hcc == _T_8[7:0] ? content_204 : _GEN_971; // @[Cat.scala 29:58]
  wire  _GEN_973 = 8'hcd == _T_8[7:0] ? content_205 : _GEN_972; // @[Cat.scala 29:58]
  wire  _GEN_974 = 8'hce == _T_8[7:0] ? content_206 : _GEN_973; // @[Cat.scala 29:58]
  wire  _GEN_975 = 8'hcf == _T_8[7:0] ? content_207 : _GEN_974; // @[Cat.scala 29:58]
  wire  _GEN_976 = 8'hd0 == _T_8[7:0] ? content_208 : _GEN_975; // @[Cat.scala 29:58]
  wire  _GEN_977 = 8'hd1 == _T_8[7:0] ? content_209 : _GEN_976; // @[Cat.scala 29:58]
  wire  _GEN_978 = 8'hd2 == _T_8[7:0] ? content_210 : _GEN_977; // @[Cat.scala 29:58]
  wire  _GEN_979 = 8'hd3 == _T_8[7:0] ? content_211 : _GEN_978; // @[Cat.scala 29:58]
  wire  _GEN_980 = 8'hd4 == _T_8[7:0] ? content_212 : _GEN_979; // @[Cat.scala 29:58]
  wire  _GEN_981 = 8'hd5 == _T_8[7:0] ? content_213 : _GEN_980; // @[Cat.scala 29:58]
  wire  _GEN_982 = 8'hd6 == _T_8[7:0] ? content_214 : _GEN_981; // @[Cat.scala 29:58]
  wire  _GEN_983 = 8'hd7 == _T_8[7:0] ? content_215 : _GEN_982; // @[Cat.scala 29:58]
  wire  _GEN_984 = 8'hd8 == _T_8[7:0] ? content_216 : _GEN_983; // @[Cat.scala 29:58]
  wire  _GEN_985 = 8'hd9 == _T_8[7:0] ? content_217 : _GEN_984; // @[Cat.scala 29:58]
  wire  _GEN_986 = 8'hda == _T_8[7:0] ? content_218 : _GEN_985; // @[Cat.scala 29:58]
  wire  _GEN_987 = 8'hdb == _T_8[7:0] ? content_219 : _GEN_986; // @[Cat.scala 29:58]
  wire  _GEN_988 = 8'hdc == _T_8[7:0] ? content_220 : _GEN_987; // @[Cat.scala 29:58]
  wire  _GEN_989 = 8'hdd == _T_8[7:0] ? content_221 : _GEN_988; // @[Cat.scala 29:58]
  wire  _GEN_990 = 8'hde == _T_8[7:0] ? content_222 : _GEN_989; // @[Cat.scala 29:58]
  wire  _GEN_991 = 8'hdf == _T_8[7:0] ? content_223 : _GEN_990; // @[Cat.scala 29:58]
  wire  _GEN_992 = 8'he0 == _T_8[7:0] ? content_224 : _GEN_991; // @[Cat.scala 29:58]
  wire  _GEN_993 = 8'he1 == _T_8[7:0] ? content_225 : _GEN_992; // @[Cat.scala 29:58]
  wire  _GEN_994 = 8'he2 == _T_8[7:0] ? content_226 : _GEN_993; // @[Cat.scala 29:58]
  wire  _GEN_995 = 8'he3 == _T_8[7:0] ? content_227 : _GEN_994; // @[Cat.scala 29:58]
  wire  _GEN_996 = 8'he4 == _T_8[7:0] ? content_228 : _GEN_995; // @[Cat.scala 29:58]
  wire  _GEN_997 = 8'he5 == _T_8[7:0] ? content_229 : _GEN_996; // @[Cat.scala 29:58]
  wire  _GEN_998 = 8'he6 == _T_8[7:0] ? content_230 : _GEN_997; // @[Cat.scala 29:58]
  wire  _GEN_999 = 8'he7 == _T_8[7:0] ? content_231 : _GEN_998; // @[Cat.scala 29:58]
  wire  _GEN_1000 = 8'he8 == _T_8[7:0] ? content_232 : _GEN_999; // @[Cat.scala 29:58]
  wire  _GEN_1001 = 8'he9 == _T_8[7:0] ? content_233 : _GEN_1000; // @[Cat.scala 29:58]
  wire  _GEN_1002 = 8'hea == _T_8[7:0] ? content_234 : _GEN_1001; // @[Cat.scala 29:58]
  wire  _GEN_1003 = 8'heb == _T_8[7:0] ? content_235 : _GEN_1002; // @[Cat.scala 29:58]
  wire  _GEN_1004 = 8'hec == _T_8[7:0] ? content_236 : _GEN_1003; // @[Cat.scala 29:58]
  wire  _GEN_1005 = 8'hed == _T_8[7:0] ? content_237 : _GEN_1004; // @[Cat.scala 29:58]
  wire  _GEN_1006 = 8'hee == _T_8[7:0] ? content_238 : _GEN_1005; // @[Cat.scala 29:58]
  wire  _GEN_1007 = 8'hef == _T_8[7:0] ? content_239 : _GEN_1006; // @[Cat.scala 29:58]
  wire  _GEN_1008 = 8'hf0 == _T_8[7:0] ? content_240 : _GEN_1007; // @[Cat.scala 29:58]
  wire  _GEN_1009 = 8'hf1 == _T_8[7:0] ? content_241 : _GEN_1008; // @[Cat.scala 29:58]
  wire  _GEN_1010 = 8'hf2 == _T_8[7:0] ? content_242 : _GEN_1009; // @[Cat.scala 29:58]
  wire  _GEN_1011 = 8'hf3 == _T_8[7:0] ? content_243 : _GEN_1010; // @[Cat.scala 29:58]
  wire  _GEN_1012 = 8'hf4 == _T_8[7:0] ? content_244 : _GEN_1011; // @[Cat.scala 29:58]
  wire  _GEN_1013 = 8'hf5 == _T_8[7:0] ? content_245 : _GEN_1012; // @[Cat.scala 29:58]
  wire  _GEN_1014 = 8'hf6 == _T_8[7:0] ? content_246 : _GEN_1013; // @[Cat.scala 29:58]
  wire  _GEN_1015 = 8'hf7 == _T_8[7:0] ? content_247 : _GEN_1014; // @[Cat.scala 29:58]
  wire  _GEN_1016 = 8'hf8 == _T_8[7:0] ? content_248 : _GEN_1015; // @[Cat.scala 29:58]
  wire  _GEN_1017 = 8'hf9 == _T_8[7:0] ? content_249 : _GEN_1016; // @[Cat.scala 29:58]
  wire  _GEN_1018 = 8'hfa == _T_8[7:0] ? content_250 : _GEN_1017; // @[Cat.scala 29:58]
  wire  _GEN_1019 = 8'hfb == _T_8[7:0] ? content_251 : _GEN_1018; // @[Cat.scala 29:58]
  wire  _GEN_1020 = 8'hfc == _T_8[7:0] ? content_252 : _GEN_1019; // @[Cat.scala 29:58]
  wire  _GEN_1021 = 8'hfd == _T_8[7:0] ? content_253 : _GEN_1020; // @[Cat.scala 29:58]
  wire  _GEN_1022 = 8'hfe == _T_8[7:0] ? content_254 : _GEN_1021; // @[Cat.scala 29:58]
  wire  _GEN_1023 = 8'hff == _T_8[7:0] ? content_255 : _GEN_1022; // @[Cat.scala 29:58]
  wire [3:0] _T_15 = {_GEN_767,_GEN_1023,_GEN_255,_GEN_511}; // @[Cat.scala 29:58]
  wire [64:0] _T_32 = {{1'd0}, io_port_1_read_in_bits_addr}; // @[elements.scala 118:104]
  wire [63:0] _T_36 = io_port_1_read_in_bits_addr + 64'h1; // @[elements.scala 118:104]
  wire [63:0] _T_39 = io_port_1_read_in_bits_addr + 64'h2; // @[elements.scala 118:104]
  wire [63:0] _T_42 = io_port_1_read_in_bits_addr + 64'h3; // @[elements.scala 118:104]
  wire  _GEN_1541 = 8'h1 == _T_36[7:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_1542 = 8'h2 == _T_36[7:0] ? content_2 : _GEN_1541; // @[Cat.scala 29:58]
  wire  _GEN_1543 = 8'h3 == _T_36[7:0] ? content_3 : _GEN_1542; // @[Cat.scala 29:58]
  wire  _GEN_1544 = 8'h4 == _T_36[7:0] ? content_4 : _GEN_1543; // @[Cat.scala 29:58]
  wire  _GEN_1545 = 8'h5 == _T_36[7:0] ? content_5 : _GEN_1544; // @[Cat.scala 29:58]
  wire  _GEN_1546 = 8'h6 == _T_36[7:0] ? content_6 : _GEN_1545; // @[Cat.scala 29:58]
  wire  _GEN_1547 = 8'h7 == _T_36[7:0] ? content_7 : _GEN_1546; // @[Cat.scala 29:58]
  wire  _GEN_1548 = 8'h8 == _T_36[7:0] ? content_8 : _GEN_1547; // @[Cat.scala 29:58]
  wire  _GEN_1549 = 8'h9 == _T_36[7:0] ? content_9 : _GEN_1548; // @[Cat.scala 29:58]
  wire  _GEN_1550 = 8'ha == _T_36[7:0] ? content_10 : _GEN_1549; // @[Cat.scala 29:58]
  wire  _GEN_1551 = 8'hb == _T_36[7:0] ? content_11 : _GEN_1550; // @[Cat.scala 29:58]
  wire  _GEN_1552 = 8'hc == _T_36[7:0] ? content_12 : _GEN_1551; // @[Cat.scala 29:58]
  wire  _GEN_1553 = 8'hd == _T_36[7:0] ? content_13 : _GEN_1552; // @[Cat.scala 29:58]
  wire  _GEN_1554 = 8'he == _T_36[7:0] ? content_14 : _GEN_1553; // @[Cat.scala 29:58]
  wire  _GEN_1555 = 8'hf == _T_36[7:0] ? content_15 : _GEN_1554; // @[Cat.scala 29:58]
  wire  _GEN_1556 = 8'h10 == _T_36[7:0] ? content_16 : _GEN_1555; // @[Cat.scala 29:58]
  wire  _GEN_1557 = 8'h11 == _T_36[7:0] ? content_17 : _GEN_1556; // @[Cat.scala 29:58]
  wire  _GEN_1558 = 8'h12 == _T_36[7:0] ? content_18 : _GEN_1557; // @[Cat.scala 29:58]
  wire  _GEN_1559 = 8'h13 == _T_36[7:0] ? content_19 : _GEN_1558; // @[Cat.scala 29:58]
  wire  _GEN_1560 = 8'h14 == _T_36[7:0] ? content_20 : _GEN_1559; // @[Cat.scala 29:58]
  wire  _GEN_1561 = 8'h15 == _T_36[7:0] ? content_21 : _GEN_1560; // @[Cat.scala 29:58]
  wire  _GEN_1562 = 8'h16 == _T_36[7:0] ? content_22 : _GEN_1561; // @[Cat.scala 29:58]
  wire  _GEN_1563 = 8'h17 == _T_36[7:0] ? content_23 : _GEN_1562; // @[Cat.scala 29:58]
  wire  _GEN_1564 = 8'h18 == _T_36[7:0] ? content_24 : _GEN_1563; // @[Cat.scala 29:58]
  wire  _GEN_1565 = 8'h19 == _T_36[7:0] ? content_25 : _GEN_1564; // @[Cat.scala 29:58]
  wire  _GEN_1566 = 8'h1a == _T_36[7:0] ? content_26 : _GEN_1565; // @[Cat.scala 29:58]
  wire  _GEN_1567 = 8'h1b == _T_36[7:0] ? content_27 : _GEN_1566; // @[Cat.scala 29:58]
  wire  _GEN_1568 = 8'h1c == _T_36[7:0] ? content_28 : _GEN_1567; // @[Cat.scala 29:58]
  wire  _GEN_1569 = 8'h1d == _T_36[7:0] ? content_29 : _GEN_1568; // @[Cat.scala 29:58]
  wire  _GEN_1570 = 8'h1e == _T_36[7:0] ? content_30 : _GEN_1569; // @[Cat.scala 29:58]
  wire  _GEN_1571 = 8'h1f == _T_36[7:0] ? content_31 : _GEN_1570; // @[Cat.scala 29:58]
  wire  _GEN_1572 = 8'h20 == _T_36[7:0] ? content_32 : _GEN_1571; // @[Cat.scala 29:58]
  wire  _GEN_1573 = 8'h21 == _T_36[7:0] ? content_33 : _GEN_1572; // @[Cat.scala 29:58]
  wire  _GEN_1574 = 8'h22 == _T_36[7:0] ? content_34 : _GEN_1573; // @[Cat.scala 29:58]
  wire  _GEN_1575 = 8'h23 == _T_36[7:0] ? content_35 : _GEN_1574; // @[Cat.scala 29:58]
  wire  _GEN_1576 = 8'h24 == _T_36[7:0] ? content_36 : _GEN_1575; // @[Cat.scala 29:58]
  wire  _GEN_1577 = 8'h25 == _T_36[7:0] ? content_37 : _GEN_1576; // @[Cat.scala 29:58]
  wire  _GEN_1578 = 8'h26 == _T_36[7:0] ? content_38 : _GEN_1577; // @[Cat.scala 29:58]
  wire  _GEN_1579 = 8'h27 == _T_36[7:0] ? content_39 : _GEN_1578; // @[Cat.scala 29:58]
  wire  _GEN_1580 = 8'h28 == _T_36[7:0] ? content_40 : _GEN_1579; // @[Cat.scala 29:58]
  wire  _GEN_1581 = 8'h29 == _T_36[7:0] ? content_41 : _GEN_1580; // @[Cat.scala 29:58]
  wire  _GEN_1582 = 8'h2a == _T_36[7:0] ? content_42 : _GEN_1581; // @[Cat.scala 29:58]
  wire  _GEN_1583 = 8'h2b == _T_36[7:0] ? content_43 : _GEN_1582; // @[Cat.scala 29:58]
  wire  _GEN_1584 = 8'h2c == _T_36[7:0] ? content_44 : _GEN_1583; // @[Cat.scala 29:58]
  wire  _GEN_1585 = 8'h2d == _T_36[7:0] ? content_45 : _GEN_1584; // @[Cat.scala 29:58]
  wire  _GEN_1586 = 8'h2e == _T_36[7:0] ? content_46 : _GEN_1585; // @[Cat.scala 29:58]
  wire  _GEN_1587 = 8'h2f == _T_36[7:0] ? content_47 : _GEN_1586; // @[Cat.scala 29:58]
  wire  _GEN_1588 = 8'h30 == _T_36[7:0] ? content_48 : _GEN_1587; // @[Cat.scala 29:58]
  wire  _GEN_1589 = 8'h31 == _T_36[7:0] ? content_49 : _GEN_1588; // @[Cat.scala 29:58]
  wire  _GEN_1590 = 8'h32 == _T_36[7:0] ? content_50 : _GEN_1589; // @[Cat.scala 29:58]
  wire  _GEN_1591 = 8'h33 == _T_36[7:0] ? content_51 : _GEN_1590; // @[Cat.scala 29:58]
  wire  _GEN_1592 = 8'h34 == _T_36[7:0] ? content_52 : _GEN_1591; // @[Cat.scala 29:58]
  wire  _GEN_1593 = 8'h35 == _T_36[7:0] ? content_53 : _GEN_1592; // @[Cat.scala 29:58]
  wire  _GEN_1594 = 8'h36 == _T_36[7:0] ? content_54 : _GEN_1593; // @[Cat.scala 29:58]
  wire  _GEN_1595 = 8'h37 == _T_36[7:0] ? content_55 : _GEN_1594; // @[Cat.scala 29:58]
  wire  _GEN_1596 = 8'h38 == _T_36[7:0] ? content_56 : _GEN_1595; // @[Cat.scala 29:58]
  wire  _GEN_1597 = 8'h39 == _T_36[7:0] ? content_57 : _GEN_1596; // @[Cat.scala 29:58]
  wire  _GEN_1598 = 8'h3a == _T_36[7:0] ? content_58 : _GEN_1597; // @[Cat.scala 29:58]
  wire  _GEN_1599 = 8'h3b == _T_36[7:0] ? content_59 : _GEN_1598; // @[Cat.scala 29:58]
  wire  _GEN_1600 = 8'h3c == _T_36[7:0] ? content_60 : _GEN_1599; // @[Cat.scala 29:58]
  wire  _GEN_1601 = 8'h3d == _T_36[7:0] ? content_61 : _GEN_1600; // @[Cat.scala 29:58]
  wire  _GEN_1602 = 8'h3e == _T_36[7:0] ? content_62 : _GEN_1601; // @[Cat.scala 29:58]
  wire  _GEN_1603 = 8'h3f == _T_36[7:0] ? content_63 : _GEN_1602; // @[Cat.scala 29:58]
  wire  _GEN_1604 = 8'h40 == _T_36[7:0] ? content_64 : _GEN_1603; // @[Cat.scala 29:58]
  wire  _GEN_1605 = 8'h41 == _T_36[7:0] ? content_65 : _GEN_1604; // @[Cat.scala 29:58]
  wire  _GEN_1606 = 8'h42 == _T_36[7:0] ? content_66 : _GEN_1605; // @[Cat.scala 29:58]
  wire  _GEN_1607 = 8'h43 == _T_36[7:0] ? content_67 : _GEN_1606; // @[Cat.scala 29:58]
  wire  _GEN_1608 = 8'h44 == _T_36[7:0] ? content_68 : _GEN_1607; // @[Cat.scala 29:58]
  wire  _GEN_1609 = 8'h45 == _T_36[7:0] ? content_69 : _GEN_1608; // @[Cat.scala 29:58]
  wire  _GEN_1610 = 8'h46 == _T_36[7:0] ? content_70 : _GEN_1609; // @[Cat.scala 29:58]
  wire  _GEN_1611 = 8'h47 == _T_36[7:0] ? content_71 : _GEN_1610; // @[Cat.scala 29:58]
  wire  _GEN_1612 = 8'h48 == _T_36[7:0] ? content_72 : _GEN_1611; // @[Cat.scala 29:58]
  wire  _GEN_1613 = 8'h49 == _T_36[7:0] ? content_73 : _GEN_1612; // @[Cat.scala 29:58]
  wire  _GEN_1614 = 8'h4a == _T_36[7:0] ? content_74 : _GEN_1613; // @[Cat.scala 29:58]
  wire  _GEN_1615 = 8'h4b == _T_36[7:0] ? content_75 : _GEN_1614; // @[Cat.scala 29:58]
  wire  _GEN_1616 = 8'h4c == _T_36[7:0] ? content_76 : _GEN_1615; // @[Cat.scala 29:58]
  wire  _GEN_1617 = 8'h4d == _T_36[7:0] ? content_77 : _GEN_1616; // @[Cat.scala 29:58]
  wire  _GEN_1618 = 8'h4e == _T_36[7:0] ? content_78 : _GEN_1617; // @[Cat.scala 29:58]
  wire  _GEN_1619 = 8'h4f == _T_36[7:0] ? content_79 : _GEN_1618; // @[Cat.scala 29:58]
  wire  _GEN_1620 = 8'h50 == _T_36[7:0] ? content_80 : _GEN_1619; // @[Cat.scala 29:58]
  wire  _GEN_1621 = 8'h51 == _T_36[7:0] ? content_81 : _GEN_1620; // @[Cat.scala 29:58]
  wire  _GEN_1622 = 8'h52 == _T_36[7:0] ? content_82 : _GEN_1621; // @[Cat.scala 29:58]
  wire  _GEN_1623 = 8'h53 == _T_36[7:0] ? content_83 : _GEN_1622; // @[Cat.scala 29:58]
  wire  _GEN_1624 = 8'h54 == _T_36[7:0] ? content_84 : _GEN_1623; // @[Cat.scala 29:58]
  wire  _GEN_1625 = 8'h55 == _T_36[7:0] ? content_85 : _GEN_1624; // @[Cat.scala 29:58]
  wire  _GEN_1626 = 8'h56 == _T_36[7:0] ? content_86 : _GEN_1625; // @[Cat.scala 29:58]
  wire  _GEN_1627 = 8'h57 == _T_36[7:0] ? content_87 : _GEN_1626; // @[Cat.scala 29:58]
  wire  _GEN_1628 = 8'h58 == _T_36[7:0] ? content_88 : _GEN_1627; // @[Cat.scala 29:58]
  wire  _GEN_1629 = 8'h59 == _T_36[7:0] ? content_89 : _GEN_1628; // @[Cat.scala 29:58]
  wire  _GEN_1630 = 8'h5a == _T_36[7:0] ? content_90 : _GEN_1629; // @[Cat.scala 29:58]
  wire  _GEN_1631 = 8'h5b == _T_36[7:0] ? content_91 : _GEN_1630; // @[Cat.scala 29:58]
  wire  _GEN_1632 = 8'h5c == _T_36[7:0] ? content_92 : _GEN_1631; // @[Cat.scala 29:58]
  wire  _GEN_1633 = 8'h5d == _T_36[7:0] ? content_93 : _GEN_1632; // @[Cat.scala 29:58]
  wire  _GEN_1634 = 8'h5e == _T_36[7:0] ? content_94 : _GEN_1633; // @[Cat.scala 29:58]
  wire  _GEN_1635 = 8'h5f == _T_36[7:0] ? content_95 : _GEN_1634; // @[Cat.scala 29:58]
  wire  _GEN_1636 = 8'h60 == _T_36[7:0] ? content_96 : _GEN_1635; // @[Cat.scala 29:58]
  wire  _GEN_1637 = 8'h61 == _T_36[7:0] ? content_97 : _GEN_1636; // @[Cat.scala 29:58]
  wire  _GEN_1638 = 8'h62 == _T_36[7:0] ? content_98 : _GEN_1637; // @[Cat.scala 29:58]
  wire  _GEN_1639 = 8'h63 == _T_36[7:0] ? content_99 : _GEN_1638; // @[Cat.scala 29:58]
  wire  _GEN_1640 = 8'h64 == _T_36[7:0] ? content_100 : _GEN_1639; // @[Cat.scala 29:58]
  wire  _GEN_1641 = 8'h65 == _T_36[7:0] ? content_101 : _GEN_1640; // @[Cat.scala 29:58]
  wire  _GEN_1642 = 8'h66 == _T_36[7:0] ? content_102 : _GEN_1641; // @[Cat.scala 29:58]
  wire  _GEN_1643 = 8'h67 == _T_36[7:0] ? content_103 : _GEN_1642; // @[Cat.scala 29:58]
  wire  _GEN_1644 = 8'h68 == _T_36[7:0] ? content_104 : _GEN_1643; // @[Cat.scala 29:58]
  wire  _GEN_1645 = 8'h69 == _T_36[7:0] ? content_105 : _GEN_1644; // @[Cat.scala 29:58]
  wire  _GEN_1646 = 8'h6a == _T_36[7:0] ? content_106 : _GEN_1645; // @[Cat.scala 29:58]
  wire  _GEN_1647 = 8'h6b == _T_36[7:0] ? content_107 : _GEN_1646; // @[Cat.scala 29:58]
  wire  _GEN_1648 = 8'h6c == _T_36[7:0] ? content_108 : _GEN_1647; // @[Cat.scala 29:58]
  wire  _GEN_1649 = 8'h6d == _T_36[7:0] ? content_109 : _GEN_1648; // @[Cat.scala 29:58]
  wire  _GEN_1650 = 8'h6e == _T_36[7:0] ? content_110 : _GEN_1649; // @[Cat.scala 29:58]
  wire  _GEN_1651 = 8'h6f == _T_36[7:0] ? content_111 : _GEN_1650; // @[Cat.scala 29:58]
  wire  _GEN_1652 = 8'h70 == _T_36[7:0] ? content_112 : _GEN_1651; // @[Cat.scala 29:58]
  wire  _GEN_1653 = 8'h71 == _T_36[7:0] ? content_113 : _GEN_1652; // @[Cat.scala 29:58]
  wire  _GEN_1654 = 8'h72 == _T_36[7:0] ? content_114 : _GEN_1653; // @[Cat.scala 29:58]
  wire  _GEN_1655 = 8'h73 == _T_36[7:0] ? content_115 : _GEN_1654; // @[Cat.scala 29:58]
  wire  _GEN_1656 = 8'h74 == _T_36[7:0] ? content_116 : _GEN_1655; // @[Cat.scala 29:58]
  wire  _GEN_1657 = 8'h75 == _T_36[7:0] ? content_117 : _GEN_1656; // @[Cat.scala 29:58]
  wire  _GEN_1658 = 8'h76 == _T_36[7:0] ? content_118 : _GEN_1657; // @[Cat.scala 29:58]
  wire  _GEN_1659 = 8'h77 == _T_36[7:0] ? content_119 : _GEN_1658; // @[Cat.scala 29:58]
  wire  _GEN_1660 = 8'h78 == _T_36[7:0] ? content_120 : _GEN_1659; // @[Cat.scala 29:58]
  wire  _GEN_1661 = 8'h79 == _T_36[7:0] ? content_121 : _GEN_1660; // @[Cat.scala 29:58]
  wire  _GEN_1662 = 8'h7a == _T_36[7:0] ? content_122 : _GEN_1661; // @[Cat.scala 29:58]
  wire  _GEN_1663 = 8'h7b == _T_36[7:0] ? content_123 : _GEN_1662; // @[Cat.scala 29:58]
  wire  _GEN_1664 = 8'h7c == _T_36[7:0] ? content_124 : _GEN_1663; // @[Cat.scala 29:58]
  wire  _GEN_1665 = 8'h7d == _T_36[7:0] ? content_125 : _GEN_1664; // @[Cat.scala 29:58]
  wire  _GEN_1666 = 8'h7e == _T_36[7:0] ? content_126 : _GEN_1665; // @[Cat.scala 29:58]
  wire  _GEN_1667 = 8'h7f == _T_36[7:0] ? content_127 : _GEN_1666; // @[Cat.scala 29:58]
  wire  _GEN_1668 = 8'h80 == _T_36[7:0] ? content_128 : _GEN_1667; // @[Cat.scala 29:58]
  wire  _GEN_1669 = 8'h81 == _T_36[7:0] ? content_129 : _GEN_1668; // @[Cat.scala 29:58]
  wire  _GEN_1670 = 8'h82 == _T_36[7:0] ? content_130 : _GEN_1669; // @[Cat.scala 29:58]
  wire  _GEN_1671 = 8'h83 == _T_36[7:0] ? content_131 : _GEN_1670; // @[Cat.scala 29:58]
  wire  _GEN_1672 = 8'h84 == _T_36[7:0] ? content_132 : _GEN_1671; // @[Cat.scala 29:58]
  wire  _GEN_1673 = 8'h85 == _T_36[7:0] ? content_133 : _GEN_1672; // @[Cat.scala 29:58]
  wire  _GEN_1674 = 8'h86 == _T_36[7:0] ? content_134 : _GEN_1673; // @[Cat.scala 29:58]
  wire  _GEN_1675 = 8'h87 == _T_36[7:0] ? content_135 : _GEN_1674; // @[Cat.scala 29:58]
  wire  _GEN_1676 = 8'h88 == _T_36[7:0] ? content_136 : _GEN_1675; // @[Cat.scala 29:58]
  wire  _GEN_1677 = 8'h89 == _T_36[7:0] ? content_137 : _GEN_1676; // @[Cat.scala 29:58]
  wire  _GEN_1678 = 8'h8a == _T_36[7:0] ? content_138 : _GEN_1677; // @[Cat.scala 29:58]
  wire  _GEN_1679 = 8'h8b == _T_36[7:0] ? content_139 : _GEN_1678; // @[Cat.scala 29:58]
  wire  _GEN_1680 = 8'h8c == _T_36[7:0] ? content_140 : _GEN_1679; // @[Cat.scala 29:58]
  wire  _GEN_1681 = 8'h8d == _T_36[7:0] ? content_141 : _GEN_1680; // @[Cat.scala 29:58]
  wire  _GEN_1682 = 8'h8e == _T_36[7:0] ? content_142 : _GEN_1681; // @[Cat.scala 29:58]
  wire  _GEN_1683 = 8'h8f == _T_36[7:0] ? content_143 : _GEN_1682; // @[Cat.scala 29:58]
  wire  _GEN_1684 = 8'h90 == _T_36[7:0] ? content_144 : _GEN_1683; // @[Cat.scala 29:58]
  wire  _GEN_1685 = 8'h91 == _T_36[7:0] ? content_145 : _GEN_1684; // @[Cat.scala 29:58]
  wire  _GEN_1686 = 8'h92 == _T_36[7:0] ? content_146 : _GEN_1685; // @[Cat.scala 29:58]
  wire  _GEN_1687 = 8'h93 == _T_36[7:0] ? content_147 : _GEN_1686; // @[Cat.scala 29:58]
  wire  _GEN_1688 = 8'h94 == _T_36[7:0] ? content_148 : _GEN_1687; // @[Cat.scala 29:58]
  wire  _GEN_1689 = 8'h95 == _T_36[7:0] ? content_149 : _GEN_1688; // @[Cat.scala 29:58]
  wire  _GEN_1690 = 8'h96 == _T_36[7:0] ? content_150 : _GEN_1689; // @[Cat.scala 29:58]
  wire  _GEN_1691 = 8'h97 == _T_36[7:0] ? content_151 : _GEN_1690; // @[Cat.scala 29:58]
  wire  _GEN_1692 = 8'h98 == _T_36[7:0] ? content_152 : _GEN_1691; // @[Cat.scala 29:58]
  wire  _GEN_1693 = 8'h99 == _T_36[7:0] ? content_153 : _GEN_1692; // @[Cat.scala 29:58]
  wire  _GEN_1694 = 8'h9a == _T_36[7:0] ? content_154 : _GEN_1693; // @[Cat.scala 29:58]
  wire  _GEN_1695 = 8'h9b == _T_36[7:0] ? content_155 : _GEN_1694; // @[Cat.scala 29:58]
  wire  _GEN_1696 = 8'h9c == _T_36[7:0] ? content_156 : _GEN_1695; // @[Cat.scala 29:58]
  wire  _GEN_1697 = 8'h9d == _T_36[7:0] ? content_157 : _GEN_1696; // @[Cat.scala 29:58]
  wire  _GEN_1698 = 8'h9e == _T_36[7:0] ? content_158 : _GEN_1697; // @[Cat.scala 29:58]
  wire  _GEN_1699 = 8'h9f == _T_36[7:0] ? content_159 : _GEN_1698; // @[Cat.scala 29:58]
  wire  _GEN_1700 = 8'ha0 == _T_36[7:0] ? content_160 : _GEN_1699; // @[Cat.scala 29:58]
  wire  _GEN_1701 = 8'ha1 == _T_36[7:0] ? content_161 : _GEN_1700; // @[Cat.scala 29:58]
  wire  _GEN_1702 = 8'ha2 == _T_36[7:0] ? content_162 : _GEN_1701; // @[Cat.scala 29:58]
  wire  _GEN_1703 = 8'ha3 == _T_36[7:0] ? content_163 : _GEN_1702; // @[Cat.scala 29:58]
  wire  _GEN_1704 = 8'ha4 == _T_36[7:0] ? content_164 : _GEN_1703; // @[Cat.scala 29:58]
  wire  _GEN_1705 = 8'ha5 == _T_36[7:0] ? content_165 : _GEN_1704; // @[Cat.scala 29:58]
  wire  _GEN_1706 = 8'ha6 == _T_36[7:0] ? content_166 : _GEN_1705; // @[Cat.scala 29:58]
  wire  _GEN_1707 = 8'ha7 == _T_36[7:0] ? content_167 : _GEN_1706; // @[Cat.scala 29:58]
  wire  _GEN_1708 = 8'ha8 == _T_36[7:0] ? content_168 : _GEN_1707; // @[Cat.scala 29:58]
  wire  _GEN_1709 = 8'ha9 == _T_36[7:0] ? content_169 : _GEN_1708; // @[Cat.scala 29:58]
  wire  _GEN_1710 = 8'haa == _T_36[7:0] ? content_170 : _GEN_1709; // @[Cat.scala 29:58]
  wire  _GEN_1711 = 8'hab == _T_36[7:0] ? content_171 : _GEN_1710; // @[Cat.scala 29:58]
  wire  _GEN_1712 = 8'hac == _T_36[7:0] ? content_172 : _GEN_1711; // @[Cat.scala 29:58]
  wire  _GEN_1713 = 8'had == _T_36[7:0] ? content_173 : _GEN_1712; // @[Cat.scala 29:58]
  wire  _GEN_1714 = 8'hae == _T_36[7:0] ? content_174 : _GEN_1713; // @[Cat.scala 29:58]
  wire  _GEN_1715 = 8'haf == _T_36[7:0] ? content_175 : _GEN_1714; // @[Cat.scala 29:58]
  wire  _GEN_1716 = 8'hb0 == _T_36[7:0] ? content_176 : _GEN_1715; // @[Cat.scala 29:58]
  wire  _GEN_1717 = 8'hb1 == _T_36[7:0] ? content_177 : _GEN_1716; // @[Cat.scala 29:58]
  wire  _GEN_1718 = 8'hb2 == _T_36[7:0] ? content_178 : _GEN_1717; // @[Cat.scala 29:58]
  wire  _GEN_1719 = 8'hb3 == _T_36[7:0] ? content_179 : _GEN_1718; // @[Cat.scala 29:58]
  wire  _GEN_1720 = 8'hb4 == _T_36[7:0] ? content_180 : _GEN_1719; // @[Cat.scala 29:58]
  wire  _GEN_1721 = 8'hb5 == _T_36[7:0] ? content_181 : _GEN_1720; // @[Cat.scala 29:58]
  wire  _GEN_1722 = 8'hb6 == _T_36[7:0] ? content_182 : _GEN_1721; // @[Cat.scala 29:58]
  wire  _GEN_1723 = 8'hb7 == _T_36[7:0] ? content_183 : _GEN_1722; // @[Cat.scala 29:58]
  wire  _GEN_1724 = 8'hb8 == _T_36[7:0] ? content_184 : _GEN_1723; // @[Cat.scala 29:58]
  wire  _GEN_1725 = 8'hb9 == _T_36[7:0] ? content_185 : _GEN_1724; // @[Cat.scala 29:58]
  wire  _GEN_1726 = 8'hba == _T_36[7:0] ? content_186 : _GEN_1725; // @[Cat.scala 29:58]
  wire  _GEN_1727 = 8'hbb == _T_36[7:0] ? content_187 : _GEN_1726; // @[Cat.scala 29:58]
  wire  _GEN_1728 = 8'hbc == _T_36[7:0] ? content_188 : _GEN_1727; // @[Cat.scala 29:58]
  wire  _GEN_1729 = 8'hbd == _T_36[7:0] ? content_189 : _GEN_1728; // @[Cat.scala 29:58]
  wire  _GEN_1730 = 8'hbe == _T_36[7:0] ? content_190 : _GEN_1729; // @[Cat.scala 29:58]
  wire  _GEN_1731 = 8'hbf == _T_36[7:0] ? content_191 : _GEN_1730; // @[Cat.scala 29:58]
  wire  _GEN_1732 = 8'hc0 == _T_36[7:0] ? content_192 : _GEN_1731; // @[Cat.scala 29:58]
  wire  _GEN_1733 = 8'hc1 == _T_36[7:0] ? content_193 : _GEN_1732; // @[Cat.scala 29:58]
  wire  _GEN_1734 = 8'hc2 == _T_36[7:0] ? content_194 : _GEN_1733; // @[Cat.scala 29:58]
  wire  _GEN_1735 = 8'hc3 == _T_36[7:0] ? content_195 : _GEN_1734; // @[Cat.scala 29:58]
  wire  _GEN_1736 = 8'hc4 == _T_36[7:0] ? content_196 : _GEN_1735; // @[Cat.scala 29:58]
  wire  _GEN_1737 = 8'hc5 == _T_36[7:0] ? content_197 : _GEN_1736; // @[Cat.scala 29:58]
  wire  _GEN_1738 = 8'hc6 == _T_36[7:0] ? content_198 : _GEN_1737; // @[Cat.scala 29:58]
  wire  _GEN_1739 = 8'hc7 == _T_36[7:0] ? content_199 : _GEN_1738; // @[Cat.scala 29:58]
  wire  _GEN_1740 = 8'hc8 == _T_36[7:0] ? content_200 : _GEN_1739; // @[Cat.scala 29:58]
  wire  _GEN_1741 = 8'hc9 == _T_36[7:0] ? content_201 : _GEN_1740; // @[Cat.scala 29:58]
  wire  _GEN_1742 = 8'hca == _T_36[7:0] ? content_202 : _GEN_1741; // @[Cat.scala 29:58]
  wire  _GEN_1743 = 8'hcb == _T_36[7:0] ? content_203 : _GEN_1742; // @[Cat.scala 29:58]
  wire  _GEN_1744 = 8'hcc == _T_36[7:0] ? content_204 : _GEN_1743; // @[Cat.scala 29:58]
  wire  _GEN_1745 = 8'hcd == _T_36[7:0] ? content_205 : _GEN_1744; // @[Cat.scala 29:58]
  wire  _GEN_1746 = 8'hce == _T_36[7:0] ? content_206 : _GEN_1745; // @[Cat.scala 29:58]
  wire  _GEN_1747 = 8'hcf == _T_36[7:0] ? content_207 : _GEN_1746; // @[Cat.scala 29:58]
  wire  _GEN_1748 = 8'hd0 == _T_36[7:0] ? content_208 : _GEN_1747; // @[Cat.scala 29:58]
  wire  _GEN_1749 = 8'hd1 == _T_36[7:0] ? content_209 : _GEN_1748; // @[Cat.scala 29:58]
  wire  _GEN_1750 = 8'hd2 == _T_36[7:0] ? content_210 : _GEN_1749; // @[Cat.scala 29:58]
  wire  _GEN_1751 = 8'hd3 == _T_36[7:0] ? content_211 : _GEN_1750; // @[Cat.scala 29:58]
  wire  _GEN_1752 = 8'hd4 == _T_36[7:0] ? content_212 : _GEN_1751; // @[Cat.scala 29:58]
  wire  _GEN_1753 = 8'hd5 == _T_36[7:0] ? content_213 : _GEN_1752; // @[Cat.scala 29:58]
  wire  _GEN_1754 = 8'hd6 == _T_36[7:0] ? content_214 : _GEN_1753; // @[Cat.scala 29:58]
  wire  _GEN_1755 = 8'hd7 == _T_36[7:0] ? content_215 : _GEN_1754; // @[Cat.scala 29:58]
  wire  _GEN_1756 = 8'hd8 == _T_36[7:0] ? content_216 : _GEN_1755; // @[Cat.scala 29:58]
  wire  _GEN_1757 = 8'hd9 == _T_36[7:0] ? content_217 : _GEN_1756; // @[Cat.scala 29:58]
  wire  _GEN_1758 = 8'hda == _T_36[7:0] ? content_218 : _GEN_1757; // @[Cat.scala 29:58]
  wire  _GEN_1759 = 8'hdb == _T_36[7:0] ? content_219 : _GEN_1758; // @[Cat.scala 29:58]
  wire  _GEN_1760 = 8'hdc == _T_36[7:0] ? content_220 : _GEN_1759; // @[Cat.scala 29:58]
  wire  _GEN_1761 = 8'hdd == _T_36[7:0] ? content_221 : _GEN_1760; // @[Cat.scala 29:58]
  wire  _GEN_1762 = 8'hde == _T_36[7:0] ? content_222 : _GEN_1761; // @[Cat.scala 29:58]
  wire  _GEN_1763 = 8'hdf == _T_36[7:0] ? content_223 : _GEN_1762; // @[Cat.scala 29:58]
  wire  _GEN_1764 = 8'he0 == _T_36[7:0] ? content_224 : _GEN_1763; // @[Cat.scala 29:58]
  wire  _GEN_1765 = 8'he1 == _T_36[7:0] ? content_225 : _GEN_1764; // @[Cat.scala 29:58]
  wire  _GEN_1766 = 8'he2 == _T_36[7:0] ? content_226 : _GEN_1765; // @[Cat.scala 29:58]
  wire  _GEN_1767 = 8'he3 == _T_36[7:0] ? content_227 : _GEN_1766; // @[Cat.scala 29:58]
  wire  _GEN_1768 = 8'he4 == _T_36[7:0] ? content_228 : _GEN_1767; // @[Cat.scala 29:58]
  wire  _GEN_1769 = 8'he5 == _T_36[7:0] ? content_229 : _GEN_1768; // @[Cat.scala 29:58]
  wire  _GEN_1770 = 8'he6 == _T_36[7:0] ? content_230 : _GEN_1769; // @[Cat.scala 29:58]
  wire  _GEN_1771 = 8'he7 == _T_36[7:0] ? content_231 : _GEN_1770; // @[Cat.scala 29:58]
  wire  _GEN_1772 = 8'he8 == _T_36[7:0] ? content_232 : _GEN_1771; // @[Cat.scala 29:58]
  wire  _GEN_1773 = 8'he9 == _T_36[7:0] ? content_233 : _GEN_1772; // @[Cat.scala 29:58]
  wire  _GEN_1774 = 8'hea == _T_36[7:0] ? content_234 : _GEN_1773; // @[Cat.scala 29:58]
  wire  _GEN_1775 = 8'heb == _T_36[7:0] ? content_235 : _GEN_1774; // @[Cat.scala 29:58]
  wire  _GEN_1776 = 8'hec == _T_36[7:0] ? content_236 : _GEN_1775; // @[Cat.scala 29:58]
  wire  _GEN_1777 = 8'hed == _T_36[7:0] ? content_237 : _GEN_1776; // @[Cat.scala 29:58]
  wire  _GEN_1778 = 8'hee == _T_36[7:0] ? content_238 : _GEN_1777; // @[Cat.scala 29:58]
  wire  _GEN_1779 = 8'hef == _T_36[7:0] ? content_239 : _GEN_1778; // @[Cat.scala 29:58]
  wire  _GEN_1780 = 8'hf0 == _T_36[7:0] ? content_240 : _GEN_1779; // @[Cat.scala 29:58]
  wire  _GEN_1781 = 8'hf1 == _T_36[7:0] ? content_241 : _GEN_1780; // @[Cat.scala 29:58]
  wire  _GEN_1782 = 8'hf2 == _T_36[7:0] ? content_242 : _GEN_1781; // @[Cat.scala 29:58]
  wire  _GEN_1783 = 8'hf3 == _T_36[7:0] ? content_243 : _GEN_1782; // @[Cat.scala 29:58]
  wire  _GEN_1784 = 8'hf4 == _T_36[7:0] ? content_244 : _GEN_1783; // @[Cat.scala 29:58]
  wire  _GEN_1785 = 8'hf5 == _T_36[7:0] ? content_245 : _GEN_1784; // @[Cat.scala 29:58]
  wire  _GEN_1786 = 8'hf6 == _T_36[7:0] ? content_246 : _GEN_1785; // @[Cat.scala 29:58]
  wire  _GEN_1787 = 8'hf7 == _T_36[7:0] ? content_247 : _GEN_1786; // @[Cat.scala 29:58]
  wire  _GEN_1788 = 8'hf8 == _T_36[7:0] ? content_248 : _GEN_1787; // @[Cat.scala 29:58]
  wire  _GEN_1789 = 8'hf9 == _T_36[7:0] ? content_249 : _GEN_1788; // @[Cat.scala 29:58]
  wire  _GEN_1790 = 8'hfa == _T_36[7:0] ? content_250 : _GEN_1789; // @[Cat.scala 29:58]
  wire  _GEN_1791 = 8'hfb == _T_36[7:0] ? content_251 : _GEN_1790; // @[Cat.scala 29:58]
  wire  _GEN_1792 = 8'hfc == _T_36[7:0] ? content_252 : _GEN_1791; // @[Cat.scala 29:58]
  wire  _GEN_1793 = 8'hfd == _T_36[7:0] ? content_253 : _GEN_1792; // @[Cat.scala 29:58]
  wire  _GEN_1794 = 8'hfe == _T_36[7:0] ? content_254 : _GEN_1793; // @[Cat.scala 29:58]
  wire  _GEN_1795 = 8'hff == _T_36[7:0] ? content_255 : _GEN_1794; // @[Cat.scala 29:58]
  wire  _GEN_1797 = 8'h1 == _T_32[7:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_1798 = 8'h2 == _T_32[7:0] ? content_2 : _GEN_1797; // @[Cat.scala 29:58]
  wire  _GEN_1799 = 8'h3 == _T_32[7:0] ? content_3 : _GEN_1798; // @[Cat.scala 29:58]
  wire  _GEN_1800 = 8'h4 == _T_32[7:0] ? content_4 : _GEN_1799; // @[Cat.scala 29:58]
  wire  _GEN_1801 = 8'h5 == _T_32[7:0] ? content_5 : _GEN_1800; // @[Cat.scala 29:58]
  wire  _GEN_1802 = 8'h6 == _T_32[7:0] ? content_6 : _GEN_1801; // @[Cat.scala 29:58]
  wire  _GEN_1803 = 8'h7 == _T_32[7:0] ? content_7 : _GEN_1802; // @[Cat.scala 29:58]
  wire  _GEN_1804 = 8'h8 == _T_32[7:0] ? content_8 : _GEN_1803; // @[Cat.scala 29:58]
  wire  _GEN_1805 = 8'h9 == _T_32[7:0] ? content_9 : _GEN_1804; // @[Cat.scala 29:58]
  wire  _GEN_1806 = 8'ha == _T_32[7:0] ? content_10 : _GEN_1805; // @[Cat.scala 29:58]
  wire  _GEN_1807 = 8'hb == _T_32[7:0] ? content_11 : _GEN_1806; // @[Cat.scala 29:58]
  wire  _GEN_1808 = 8'hc == _T_32[7:0] ? content_12 : _GEN_1807; // @[Cat.scala 29:58]
  wire  _GEN_1809 = 8'hd == _T_32[7:0] ? content_13 : _GEN_1808; // @[Cat.scala 29:58]
  wire  _GEN_1810 = 8'he == _T_32[7:0] ? content_14 : _GEN_1809; // @[Cat.scala 29:58]
  wire  _GEN_1811 = 8'hf == _T_32[7:0] ? content_15 : _GEN_1810; // @[Cat.scala 29:58]
  wire  _GEN_1812 = 8'h10 == _T_32[7:0] ? content_16 : _GEN_1811; // @[Cat.scala 29:58]
  wire  _GEN_1813 = 8'h11 == _T_32[7:0] ? content_17 : _GEN_1812; // @[Cat.scala 29:58]
  wire  _GEN_1814 = 8'h12 == _T_32[7:0] ? content_18 : _GEN_1813; // @[Cat.scala 29:58]
  wire  _GEN_1815 = 8'h13 == _T_32[7:0] ? content_19 : _GEN_1814; // @[Cat.scala 29:58]
  wire  _GEN_1816 = 8'h14 == _T_32[7:0] ? content_20 : _GEN_1815; // @[Cat.scala 29:58]
  wire  _GEN_1817 = 8'h15 == _T_32[7:0] ? content_21 : _GEN_1816; // @[Cat.scala 29:58]
  wire  _GEN_1818 = 8'h16 == _T_32[7:0] ? content_22 : _GEN_1817; // @[Cat.scala 29:58]
  wire  _GEN_1819 = 8'h17 == _T_32[7:0] ? content_23 : _GEN_1818; // @[Cat.scala 29:58]
  wire  _GEN_1820 = 8'h18 == _T_32[7:0] ? content_24 : _GEN_1819; // @[Cat.scala 29:58]
  wire  _GEN_1821 = 8'h19 == _T_32[7:0] ? content_25 : _GEN_1820; // @[Cat.scala 29:58]
  wire  _GEN_1822 = 8'h1a == _T_32[7:0] ? content_26 : _GEN_1821; // @[Cat.scala 29:58]
  wire  _GEN_1823 = 8'h1b == _T_32[7:0] ? content_27 : _GEN_1822; // @[Cat.scala 29:58]
  wire  _GEN_1824 = 8'h1c == _T_32[7:0] ? content_28 : _GEN_1823; // @[Cat.scala 29:58]
  wire  _GEN_1825 = 8'h1d == _T_32[7:0] ? content_29 : _GEN_1824; // @[Cat.scala 29:58]
  wire  _GEN_1826 = 8'h1e == _T_32[7:0] ? content_30 : _GEN_1825; // @[Cat.scala 29:58]
  wire  _GEN_1827 = 8'h1f == _T_32[7:0] ? content_31 : _GEN_1826; // @[Cat.scala 29:58]
  wire  _GEN_1828 = 8'h20 == _T_32[7:0] ? content_32 : _GEN_1827; // @[Cat.scala 29:58]
  wire  _GEN_1829 = 8'h21 == _T_32[7:0] ? content_33 : _GEN_1828; // @[Cat.scala 29:58]
  wire  _GEN_1830 = 8'h22 == _T_32[7:0] ? content_34 : _GEN_1829; // @[Cat.scala 29:58]
  wire  _GEN_1831 = 8'h23 == _T_32[7:0] ? content_35 : _GEN_1830; // @[Cat.scala 29:58]
  wire  _GEN_1832 = 8'h24 == _T_32[7:0] ? content_36 : _GEN_1831; // @[Cat.scala 29:58]
  wire  _GEN_1833 = 8'h25 == _T_32[7:0] ? content_37 : _GEN_1832; // @[Cat.scala 29:58]
  wire  _GEN_1834 = 8'h26 == _T_32[7:0] ? content_38 : _GEN_1833; // @[Cat.scala 29:58]
  wire  _GEN_1835 = 8'h27 == _T_32[7:0] ? content_39 : _GEN_1834; // @[Cat.scala 29:58]
  wire  _GEN_1836 = 8'h28 == _T_32[7:0] ? content_40 : _GEN_1835; // @[Cat.scala 29:58]
  wire  _GEN_1837 = 8'h29 == _T_32[7:0] ? content_41 : _GEN_1836; // @[Cat.scala 29:58]
  wire  _GEN_1838 = 8'h2a == _T_32[7:0] ? content_42 : _GEN_1837; // @[Cat.scala 29:58]
  wire  _GEN_1839 = 8'h2b == _T_32[7:0] ? content_43 : _GEN_1838; // @[Cat.scala 29:58]
  wire  _GEN_1840 = 8'h2c == _T_32[7:0] ? content_44 : _GEN_1839; // @[Cat.scala 29:58]
  wire  _GEN_1841 = 8'h2d == _T_32[7:0] ? content_45 : _GEN_1840; // @[Cat.scala 29:58]
  wire  _GEN_1842 = 8'h2e == _T_32[7:0] ? content_46 : _GEN_1841; // @[Cat.scala 29:58]
  wire  _GEN_1843 = 8'h2f == _T_32[7:0] ? content_47 : _GEN_1842; // @[Cat.scala 29:58]
  wire  _GEN_1844 = 8'h30 == _T_32[7:0] ? content_48 : _GEN_1843; // @[Cat.scala 29:58]
  wire  _GEN_1845 = 8'h31 == _T_32[7:0] ? content_49 : _GEN_1844; // @[Cat.scala 29:58]
  wire  _GEN_1846 = 8'h32 == _T_32[7:0] ? content_50 : _GEN_1845; // @[Cat.scala 29:58]
  wire  _GEN_1847 = 8'h33 == _T_32[7:0] ? content_51 : _GEN_1846; // @[Cat.scala 29:58]
  wire  _GEN_1848 = 8'h34 == _T_32[7:0] ? content_52 : _GEN_1847; // @[Cat.scala 29:58]
  wire  _GEN_1849 = 8'h35 == _T_32[7:0] ? content_53 : _GEN_1848; // @[Cat.scala 29:58]
  wire  _GEN_1850 = 8'h36 == _T_32[7:0] ? content_54 : _GEN_1849; // @[Cat.scala 29:58]
  wire  _GEN_1851 = 8'h37 == _T_32[7:0] ? content_55 : _GEN_1850; // @[Cat.scala 29:58]
  wire  _GEN_1852 = 8'h38 == _T_32[7:0] ? content_56 : _GEN_1851; // @[Cat.scala 29:58]
  wire  _GEN_1853 = 8'h39 == _T_32[7:0] ? content_57 : _GEN_1852; // @[Cat.scala 29:58]
  wire  _GEN_1854 = 8'h3a == _T_32[7:0] ? content_58 : _GEN_1853; // @[Cat.scala 29:58]
  wire  _GEN_1855 = 8'h3b == _T_32[7:0] ? content_59 : _GEN_1854; // @[Cat.scala 29:58]
  wire  _GEN_1856 = 8'h3c == _T_32[7:0] ? content_60 : _GEN_1855; // @[Cat.scala 29:58]
  wire  _GEN_1857 = 8'h3d == _T_32[7:0] ? content_61 : _GEN_1856; // @[Cat.scala 29:58]
  wire  _GEN_1858 = 8'h3e == _T_32[7:0] ? content_62 : _GEN_1857; // @[Cat.scala 29:58]
  wire  _GEN_1859 = 8'h3f == _T_32[7:0] ? content_63 : _GEN_1858; // @[Cat.scala 29:58]
  wire  _GEN_1860 = 8'h40 == _T_32[7:0] ? content_64 : _GEN_1859; // @[Cat.scala 29:58]
  wire  _GEN_1861 = 8'h41 == _T_32[7:0] ? content_65 : _GEN_1860; // @[Cat.scala 29:58]
  wire  _GEN_1862 = 8'h42 == _T_32[7:0] ? content_66 : _GEN_1861; // @[Cat.scala 29:58]
  wire  _GEN_1863 = 8'h43 == _T_32[7:0] ? content_67 : _GEN_1862; // @[Cat.scala 29:58]
  wire  _GEN_1864 = 8'h44 == _T_32[7:0] ? content_68 : _GEN_1863; // @[Cat.scala 29:58]
  wire  _GEN_1865 = 8'h45 == _T_32[7:0] ? content_69 : _GEN_1864; // @[Cat.scala 29:58]
  wire  _GEN_1866 = 8'h46 == _T_32[7:0] ? content_70 : _GEN_1865; // @[Cat.scala 29:58]
  wire  _GEN_1867 = 8'h47 == _T_32[7:0] ? content_71 : _GEN_1866; // @[Cat.scala 29:58]
  wire  _GEN_1868 = 8'h48 == _T_32[7:0] ? content_72 : _GEN_1867; // @[Cat.scala 29:58]
  wire  _GEN_1869 = 8'h49 == _T_32[7:0] ? content_73 : _GEN_1868; // @[Cat.scala 29:58]
  wire  _GEN_1870 = 8'h4a == _T_32[7:0] ? content_74 : _GEN_1869; // @[Cat.scala 29:58]
  wire  _GEN_1871 = 8'h4b == _T_32[7:0] ? content_75 : _GEN_1870; // @[Cat.scala 29:58]
  wire  _GEN_1872 = 8'h4c == _T_32[7:0] ? content_76 : _GEN_1871; // @[Cat.scala 29:58]
  wire  _GEN_1873 = 8'h4d == _T_32[7:0] ? content_77 : _GEN_1872; // @[Cat.scala 29:58]
  wire  _GEN_1874 = 8'h4e == _T_32[7:0] ? content_78 : _GEN_1873; // @[Cat.scala 29:58]
  wire  _GEN_1875 = 8'h4f == _T_32[7:0] ? content_79 : _GEN_1874; // @[Cat.scala 29:58]
  wire  _GEN_1876 = 8'h50 == _T_32[7:0] ? content_80 : _GEN_1875; // @[Cat.scala 29:58]
  wire  _GEN_1877 = 8'h51 == _T_32[7:0] ? content_81 : _GEN_1876; // @[Cat.scala 29:58]
  wire  _GEN_1878 = 8'h52 == _T_32[7:0] ? content_82 : _GEN_1877; // @[Cat.scala 29:58]
  wire  _GEN_1879 = 8'h53 == _T_32[7:0] ? content_83 : _GEN_1878; // @[Cat.scala 29:58]
  wire  _GEN_1880 = 8'h54 == _T_32[7:0] ? content_84 : _GEN_1879; // @[Cat.scala 29:58]
  wire  _GEN_1881 = 8'h55 == _T_32[7:0] ? content_85 : _GEN_1880; // @[Cat.scala 29:58]
  wire  _GEN_1882 = 8'h56 == _T_32[7:0] ? content_86 : _GEN_1881; // @[Cat.scala 29:58]
  wire  _GEN_1883 = 8'h57 == _T_32[7:0] ? content_87 : _GEN_1882; // @[Cat.scala 29:58]
  wire  _GEN_1884 = 8'h58 == _T_32[7:0] ? content_88 : _GEN_1883; // @[Cat.scala 29:58]
  wire  _GEN_1885 = 8'h59 == _T_32[7:0] ? content_89 : _GEN_1884; // @[Cat.scala 29:58]
  wire  _GEN_1886 = 8'h5a == _T_32[7:0] ? content_90 : _GEN_1885; // @[Cat.scala 29:58]
  wire  _GEN_1887 = 8'h5b == _T_32[7:0] ? content_91 : _GEN_1886; // @[Cat.scala 29:58]
  wire  _GEN_1888 = 8'h5c == _T_32[7:0] ? content_92 : _GEN_1887; // @[Cat.scala 29:58]
  wire  _GEN_1889 = 8'h5d == _T_32[7:0] ? content_93 : _GEN_1888; // @[Cat.scala 29:58]
  wire  _GEN_1890 = 8'h5e == _T_32[7:0] ? content_94 : _GEN_1889; // @[Cat.scala 29:58]
  wire  _GEN_1891 = 8'h5f == _T_32[7:0] ? content_95 : _GEN_1890; // @[Cat.scala 29:58]
  wire  _GEN_1892 = 8'h60 == _T_32[7:0] ? content_96 : _GEN_1891; // @[Cat.scala 29:58]
  wire  _GEN_1893 = 8'h61 == _T_32[7:0] ? content_97 : _GEN_1892; // @[Cat.scala 29:58]
  wire  _GEN_1894 = 8'h62 == _T_32[7:0] ? content_98 : _GEN_1893; // @[Cat.scala 29:58]
  wire  _GEN_1895 = 8'h63 == _T_32[7:0] ? content_99 : _GEN_1894; // @[Cat.scala 29:58]
  wire  _GEN_1896 = 8'h64 == _T_32[7:0] ? content_100 : _GEN_1895; // @[Cat.scala 29:58]
  wire  _GEN_1897 = 8'h65 == _T_32[7:0] ? content_101 : _GEN_1896; // @[Cat.scala 29:58]
  wire  _GEN_1898 = 8'h66 == _T_32[7:0] ? content_102 : _GEN_1897; // @[Cat.scala 29:58]
  wire  _GEN_1899 = 8'h67 == _T_32[7:0] ? content_103 : _GEN_1898; // @[Cat.scala 29:58]
  wire  _GEN_1900 = 8'h68 == _T_32[7:0] ? content_104 : _GEN_1899; // @[Cat.scala 29:58]
  wire  _GEN_1901 = 8'h69 == _T_32[7:0] ? content_105 : _GEN_1900; // @[Cat.scala 29:58]
  wire  _GEN_1902 = 8'h6a == _T_32[7:0] ? content_106 : _GEN_1901; // @[Cat.scala 29:58]
  wire  _GEN_1903 = 8'h6b == _T_32[7:0] ? content_107 : _GEN_1902; // @[Cat.scala 29:58]
  wire  _GEN_1904 = 8'h6c == _T_32[7:0] ? content_108 : _GEN_1903; // @[Cat.scala 29:58]
  wire  _GEN_1905 = 8'h6d == _T_32[7:0] ? content_109 : _GEN_1904; // @[Cat.scala 29:58]
  wire  _GEN_1906 = 8'h6e == _T_32[7:0] ? content_110 : _GEN_1905; // @[Cat.scala 29:58]
  wire  _GEN_1907 = 8'h6f == _T_32[7:0] ? content_111 : _GEN_1906; // @[Cat.scala 29:58]
  wire  _GEN_1908 = 8'h70 == _T_32[7:0] ? content_112 : _GEN_1907; // @[Cat.scala 29:58]
  wire  _GEN_1909 = 8'h71 == _T_32[7:0] ? content_113 : _GEN_1908; // @[Cat.scala 29:58]
  wire  _GEN_1910 = 8'h72 == _T_32[7:0] ? content_114 : _GEN_1909; // @[Cat.scala 29:58]
  wire  _GEN_1911 = 8'h73 == _T_32[7:0] ? content_115 : _GEN_1910; // @[Cat.scala 29:58]
  wire  _GEN_1912 = 8'h74 == _T_32[7:0] ? content_116 : _GEN_1911; // @[Cat.scala 29:58]
  wire  _GEN_1913 = 8'h75 == _T_32[7:0] ? content_117 : _GEN_1912; // @[Cat.scala 29:58]
  wire  _GEN_1914 = 8'h76 == _T_32[7:0] ? content_118 : _GEN_1913; // @[Cat.scala 29:58]
  wire  _GEN_1915 = 8'h77 == _T_32[7:0] ? content_119 : _GEN_1914; // @[Cat.scala 29:58]
  wire  _GEN_1916 = 8'h78 == _T_32[7:0] ? content_120 : _GEN_1915; // @[Cat.scala 29:58]
  wire  _GEN_1917 = 8'h79 == _T_32[7:0] ? content_121 : _GEN_1916; // @[Cat.scala 29:58]
  wire  _GEN_1918 = 8'h7a == _T_32[7:0] ? content_122 : _GEN_1917; // @[Cat.scala 29:58]
  wire  _GEN_1919 = 8'h7b == _T_32[7:0] ? content_123 : _GEN_1918; // @[Cat.scala 29:58]
  wire  _GEN_1920 = 8'h7c == _T_32[7:0] ? content_124 : _GEN_1919; // @[Cat.scala 29:58]
  wire  _GEN_1921 = 8'h7d == _T_32[7:0] ? content_125 : _GEN_1920; // @[Cat.scala 29:58]
  wire  _GEN_1922 = 8'h7e == _T_32[7:0] ? content_126 : _GEN_1921; // @[Cat.scala 29:58]
  wire  _GEN_1923 = 8'h7f == _T_32[7:0] ? content_127 : _GEN_1922; // @[Cat.scala 29:58]
  wire  _GEN_1924 = 8'h80 == _T_32[7:0] ? content_128 : _GEN_1923; // @[Cat.scala 29:58]
  wire  _GEN_1925 = 8'h81 == _T_32[7:0] ? content_129 : _GEN_1924; // @[Cat.scala 29:58]
  wire  _GEN_1926 = 8'h82 == _T_32[7:0] ? content_130 : _GEN_1925; // @[Cat.scala 29:58]
  wire  _GEN_1927 = 8'h83 == _T_32[7:0] ? content_131 : _GEN_1926; // @[Cat.scala 29:58]
  wire  _GEN_1928 = 8'h84 == _T_32[7:0] ? content_132 : _GEN_1927; // @[Cat.scala 29:58]
  wire  _GEN_1929 = 8'h85 == _T_32[7:0] ? content_133 : _GEN_1928; // @[Cat.scala 29:58]
  wire  _GEN_1930 = 8'h86 == _T_32[7:0] ? content_134 : _GEN_1929; // @[Cat.scala 29:58]
  wire  _GEN_1931 = 8'h87 == _T_32[7:0] ? content_135 : _GEN_1930; // @[Cat.scala 29:58]
  wire  _GEN_1932 = 8'h88 == _T_32[7:0] ? content_136 : _GEN_1931; // @[Cat.scala 29:58]
  wire  _GEN_1933 = 8'h89 == _T_32[7:0] ? content_137 : _GEN_1932; // @[Cat.scala 29:58]
  wire  _GEN_1934 = 8'h8a == _T_32[7:0] ? content_138 : _GEN_1933; // @[Cat.scala 29:58]
  wire  _GEN_1935 = 8'h8b == _T_32[7:0] ? content_139 : _GEN_1934; // @[Cat.scala 29:58]
  wire  _GEN_1936 = 8'h8c == _T_32[7:0] ? content_140 : _GEN_1935; // @[Cat.scala 29:58]
  wire  _GEN_1937 = 8'h8d == _T_32[7:0] ? content_141 : _GEN_1936; // @[Cat.scala 29:58]
  wire  _GEN_1938 = 8'h8e == _T_32[7:0] ? content_142 : _GEN_1937; // @[Cat.scala 29:58]
  wire  _GEN_1939 = 8'h8f == _T_32[7:0] ? content_143 : _GEN_1938; // @[Cat.scala 29:58]
  wire  _GEN_1940 = 8'h90 == _T_32[7:0] ? content_144 : _GEN_1939; // @[Cat.scala 29:58]
  wire  _GEN_1941 = 8'h91 == _T_32[7:0] ? content_145 : _GEN_1940; // @[Cat.scala 29:58]
  wire  _GEN_1942 = 8'h92 == _T_32[7:0] ? content_146 : _GEN_1941; // @[Cat.scala 29:58]
  wire  _GEN_1943 = 8'h93 == _T_32[7:0] ? content_147 : _GEN_1942; // @[Cat.scala 29:58]
  wire  _GEN_1944 = 8'h94 == _T_32[7:0] ? content_148 : _GEN_1943; // @[Cat.scala 29:58]
  wire  _GEN_1945 = 8'h95 == _T_32[7:0] ? content_149 : _GEN_1944; // @[Cat.scala 29:58]
  wire  _GEN_1946 = 8'h96 == _T_32[7:0] ? content_150 : _GEN_1945; // @[Cat.scala 29:58]
  wire  _GEN_1947 = 8'h97 == _T_32[7:0] ? content_151 : _GEN_1946; // @[Cat.scala 29:58]
  wire  _GEN_1948 = 8'h98 == _T_32[7:0] ? content_152 : _GEN_1947; // @[Cat.scala 29:58]
  wire  _GEN_1949 = 8'h99 == _T_32[7:0] ? content_153 : _GEN_1948; // @[Cat.scala 29:58]
  wire  _GEN_1950 = 8'h9a == _T_32[7:0] ? content_154 : _GEN_1949; // @[Cat.scala 29:58]
  wire  _GEN_1951 = 8'h9b == _T_32[7:0] ? content_155 : _GEN_1950; // @[Cat.scala 29:58]
  wire  _GEN_1952 = 8'h9c == _T_32[7:0] ? content_156 : _GEN_1951; // @[Cat.scala 29:58]
  wire  _GEN_1953 = 8'h9d == _T_32[7:0] ? content_157 : _GEN_1952; // @[Cat.scala 29:58]
  wire  _GEN_1954 = 8'h9e == _T_32[7:0] ? content_158 : _GEN_1953; // @[Cat.scala 29:58]
  wire  _GEN_1955 = 8'h9f == _T_32[7:0] ? content_159 : _GEN_1954; // @[Cat.scala 29:58]
  wire  _GEN_1956 = 8'ha0 == _T_32[7:0] ? content_160 : _GEN_1955; // @[Cat.scala 29:58]
  wire  _GEN_1957 = 8'ha1 == _T_32[7:0] ? content_161 : _GEN_1956; // @[Cat.scala 29:58]
  wire  _GEN_1958 = 8'ha2 == _T_32[7:0] ? content_162 : _GEN_1957; // @[Cat.scala 29:58]
  wire  _GEN_1959 = 8'ha3 == _T_32[7:0] ? content_163 : _GEN_1958; // @[Cat.scala 29:58]
  wire  _GEN_1960 = 8'ha4 == _T_32[7:0] ? content_164 : _GEN_1959; // @[Cat.scala 29:58]
  wire  _GEN_1961 = 8'ha5 == _T_32[7:0] ? content_165 : _GEN_1960; // @[Cat.scala 29:58]
  wire  _GEN_1962 = 8'ha6 == _T_32[7:0] ? content_166 : _GEN_1961; // @[Cat.scala 29:58]
  wire  _GEN_1963 = 8'ha7 == _T_32[7:0] ? content_167 : _GEN_1962; // @[Cat.scala 29:58]
  wire  _GEN_1964 = 8'ha8 == _T_32[7:0] ? content_168 : _GEN_1963; // @[Cat.scala 29:58]
  wire  _GEN_1965 = 8'ha9 == _T_32[7:0] ? content_169 : _GEN_1964; // @[Cat.scala 29:58]
  wire  _GEN_1966 = 8'haa == _T_32[7:0] ? content_170 : _GEN_1965; // @[Cat.scala 29:58]
  wire  _GEN_1967 = 8'hab == _T_32[7:0] ? content_171 : _GEN_1966; // @[Cat.scala 29:58]
  wire  _GEN_1968 = 8'hac == _T_32[7:0] ? content_172 : _GEN_1967; // @[Cat.scala 29:58]
  wire  _GEN_1969 = 8'had == _T_32[7:0] ? content_173 : _GEN_1968; // @[Cat.scala 29:58]
  wire  _GEN_1970 = 8'hae == _T_32[7:0] ? content_174 : _GEN_1969; // @[Cat.scala 29:58]
  wire  _GEN_1971 = 8'haf == _T_32[7:0] ? content_175 : _GEN_1970; // @[Cat.scala 29:58]
  wire  _GEN_1972 = 8'hb0 == _T_32[7:0] ? content_176 : _GEN_1971; // @[Cat.scala 29:58]
  wire  _GEN_1973 = 8'hb1 == _T_32[7:0] ? content_177 : _GEN_1972; // @[Cat.scala 29:58]
  wire  _GEN_1974 = 8'hb2 == _T_32[7:0] ? content_178 : _GEN_1973; // @[Cat.scala 29:58]
  wire  _GEN_1975 = 8'hb3 == _T_32[7:0] ? content_179 : _GEN_1974; // @[Cat.scala 29:58]
  wire  _GEN_1976 = 8'hb4 == _T_32[7:0] ? content_180 : _GEN_1975; // @[Cat.scala 29:58]
  wire  _GEN_1977 = 8'hb5 == _T_32[7:0] ? content_181 : _GEN_1976; // @[Cat.scala 29:58]
  wire  _GEN_1978 = 8'hb6 == _T_32[7:0] ? content_182 : _GEN_1977; // @[Cat.scala 29:58]
  wire  _GEN_1979 = 8'hb7 == _T_32[7:0] ? content_183 : _GEN_1978; // @[Cat.scala 29:58]
  wire  _GEN_1980 = 8'hb8 == _T_32[7:0] ? content_184 : _GEN_1979; // @[Cat.scala 29:58]
  wire  _GEN_1981 = 8'hb9 == _T_32[7:0] ? content_185 : _GEN_1980; // @[Cat.scala 29:58]
  wire  _GEN_1982 = 8'hba == _T_32[7:0] ? content_186 : _GEN_1981; // @[Cat.scala 29:58]
  wire  _GEN_1983 = 8'hbb == _T_32[7:0] ? content_187 : _GEN_1982; // @[Cat.scala 29:58]
  wire  _GEN_1984 = 8'hbc == _T_32[7:0] ? content_188 : _GEN_1983; // @[Cat.scala 29:58]
  wire  _GEN_1985 = 8'hbd == _T_32[7:0] ? content_189 : _GEN_1984; // @[Cat.scala 29:58]
  wire  _GEN_1986 = 8'hbe == _T_32[7:0] ? content_190 : _GEN_1985; // @[Cat.scala 29:58]
  wire  _GEN_1987 = 8'hbf == _T_32[7:0] ? content_191 : _GEN_1986; // @[Cat.scala 29:58]
  wire  _GEN_1988 = 8'hc0 == _T_32[7:0] ? content_192 : _GEN_1987; // @[Cat.scala 29:58]
  wire  _GEN_1989 = 8'hc1 == _T_32[7:0] ? content_193 : _GEN_1988; // @[Cat.scala 29:58]
  wire  _GEN_1990 = 8'hc2 == _T_32[7:0] ? content_194 : _GEN_1989; // @[Cat.scala 29:58]
  wire  _GEN_1991 = 8'hc3 == _T_32[7:0] ? content_195 : _GEN_1990; // @[Cat.scala 29:58]
  wire  _GEN_1992 = 8'hc4 == _T_32[7:0] ? content_196 : _GEN_1991; // @[Cat.scala 29:58]
  wire  _GEN_1993 = 8'hc5 == _T_32[7:0] ? content_197 : _GEN_1992; // @[Cat.scala 29:58]
  wire  _GEN_1994 = 8'hc6 == _T_32[7:0] ? content_198 : _GEN_1993; // @[Cat.scala 29:58]
  wire  _GEN_1995 = 8'hc7 == _T_32[7:0] ? content_199 : _GEN_1994; // @[Cat.scala 29:58]
  wire  _GEN_1996 = 8'hc8 == _T_32[7:0] ? content_200 : _GEN_1995; // @[Cat.scala 29:58]
  wire  _GEN_1997 = 8'hc9 == _T_32[7:0] ? content_201 : _GEN_1996; // @[Cat.scala 29:58]
  wire  _GEN_1998 = 8'hca == _T_32[7:0] ? content_202 : _GEN_1997; // @[Cat.scala 29:58]
  wire  _GEN_1999 = 8'hcb == _T_32[7:0] ? content_203 : _GEN_1998; // @[Cat.scala 29:58]
  wire  _GEN_2000 = 8'hcc == _T_32[7:0] ? content_204 : _GEN_1999; // @[Cat.scala 29:58]
  wire  _GEN_2001 = 8'hcd == _T_32[7:0] ? content_205 : _GEN_2000; // @[Cat.scala 29:58]
  wire  _GEN_2002 = 8'hce == _T_32[7:0] ? content_206 : _GEN_2001; // @[Cat.scala 29:58]
  wire  _GEN_2003 = 8'hcf == _T_32[7:0] ? content_207 : _GEN_2002; // @[Cat.scala 29:58]
  wire  _GEN_2004 = 8'hd0 == _T_32[7:0] ? content_208 : _GEN_2003; // @[Cat.scala 29:58]
  wire  _GEN_2005 = 8'hd1 == _T_32[7:0] ? content_209 : _GEN_2004; // @[Cat.scala 29:58]
  wire  _GEN_2006 = 8'hd2 == _T_32[7:0] ? content_210 : _GEN_2005; // @[Cat.scala 29:58]
  wire  _GEN_2007 = 8'hd3 == _T_32[7:0] ? content_211 : _GEN_2006; // @[Cat.scala 29:58]
  wire  _GEN_2008 = 8'hd4 == _T_32[7:0] ? content_212 : _GEN_2007; // @[Cat.scala 29:58]
  wire  _GEN_2009 = 8'hd5 == _T_32[7:0] ? content_213 : _GEN_2008; // @[Cat.scala 29:58]
  wire  _GEN_2010 = 8'hd6 == _T_32[7:0] ? content_214 : _GEN_2009; // @[Cat.scala 29:58]
  wire  _GEN_2011 = 8'hd7 == _T_32[7:0] ? content_215 : _GEN_2010; // @[Cat.scala 29:58]
  wire  _GEN_2012 = 8'hd8 == _T_32[7:0] ? content_216 : _GEN_2011; // @[Cat.scala 29:58]
  wire  _GEN_2013 = 8'hd9 == _T_32[7:0] ? content_217 : _GEN_2012; // @[Cat.scala 29:58]
  wire  _GEN_2014 = 8'hda == _T_32[7:0] ? content_218 : _GEN_2013; // @[Cat.scala 29:58]
  wire  _GEN_2015 = 8'hdb == _T_32[7:0] ? content_219 : _GEN_2014; // @[Cat.scala 29:58]
  wire  _GEN_2016 = 8'hdc == _T_32[7:0] ? content_220 : _GEN_2015; // @[Cat.scala 29:58]
  wire  _GEN_2017 = 8'hdd == _T_32[7:0] ? content_221 : _GEN_2016; // @[Cat.scala 29:58]
  wire  _GEN_2018 = 8'hde == _T_32[7:0] ? content_222 : _GEN_2017; // @[Cat.scala 29:58]
  wire  _GEN_2019 = 8'hdf == _T_32[7:0] ? content_223 : _GEN_2018; // @[Cat.scala 29:58]
  wire  _GEN_2020 = 8'he0 == _T_32[7:0] ? content_224 : _GEN_2019; // @[Cat.scala 29:58]
  wire  _GEN_2021 = 8'he1 == _T_32[7:0] ? content_225 : _GEN_2020; // @[Cat.scala 29:58]
  wire  _GEN_2022 = 8'he2 == _T_32[7:0] ? content_226 : _GEN_2021; // @[Cat.scala 29:58]
  wire  _GEN_2023 = 8'he3 == _T_32[7:0] ? content_227 : _GEN_2022; // @[Cat.scala 29:58]
  wire  _GEN_2024 = 8'he4 == _T_32[7:0] ? content_228 : _GEN_2023; // @[Cat.scala 29:58]
  wire  _GEN_2025 = 8'he5 == _T_32[7:0] ? content_229 : _GEN_2024; // @[Cat.scala 29:58]
  wire  _GEN_2026 = 8'he6 == _T_32[7:0] ? content_230 : _GEN_2025; // @[Cat.scala 29:58]
  wire  _GEN_2027 = 8'he7 == _T_32[7:0] ? content_231 : _GEN_2026; // @[Cat.scala 29:58]
  wire  _GEN_2028 = 8'he8 == _T_32[7:0] ? content_232 : _GEN_2027; // @[Cat.scala 29:58]
  wire  _GEN_2029 = 8'he9 == _T_32[7:0] ? content_233 : _GEN_2028; // @[Cat.scala 29:58]
  wire  _GEN_2030 = 8'hea == _T_32[7:0] ? content_234 : _GEN_2029; // @[Cat.scala 29:58]
  wire  _GEN_2031 = 8'heb == _T_32[7:0] ? content_235 : _GEN_2030; // @[Cat.scala 29:58]
  wire  _GEN_2032 = 8'hec == _T_32[7:0] ? content_236 : _GEN_2031; // @[Cat.scala 29:58]
  wire  _GEN_2033 = 8'hed == _T_32[7:0] ? content_237 : _GEN_2032; // @[Cat.scala 29:58]
  wire  _GEN_2034 = 8'hee == _T_32[7:0] ? content_238 : _GEN_2033; // @[Cat.scala 29:58]
  wire  _GEN_2035 = 8'hef == _T_32[7:0] ? content_239 : _GEN_2034; // @[Cat.scala 29:58]
  wire  _GEN_2036 = 8'hf0 == _T_32[7:0] ? content_240 : _GEN_2035; // @[Cat.scala 29:58]
  wire  _GEN_2037 = 8'hf1 == _T_32[7:0] ? content_241 : _GEN_2036; // @[Cat.scala 29:58]
  wire  _GEN_2038 = 8'hf2 == _T_32[7:0] ? content_242 : _GEN_2037; // @[Cat.scala 29:58]
  wire  _GEN_2039 = 8'hf3 == _T_32[7:0] ? content_243 : _GEN_2038; // @[Cat.scala 29:58]
  wire  _GEN_2040 = 8'hf4 == _T_32[7:0] ? content_244 : _GEN_2039; // @[Cat.scala 29:58]
  wire  _GEN_2041 = 8'hf5 == _T_32[7:0] ? content_245 : _GEN_2040; // @[Cat.scala 29:58]
  wire  _GEN_2042 = 8'hf6 == _T_32[7:0] ? content_246 : _GEN_2041; // @[Cat.scala 29:58]
  wire  _GEN_2043 = 8'hf7 == _T_32[7:0] ? content_247 : _GEN_2042; // @[Cat.scala 29:58]
  wire  _GEN_2044 = 8'hf8 == _T_32[7:0] ? content_248 : _GEN_2043; // @[Cat.scala 29:58]
  wire  _GEN_2045 = 8'hf9 == _T_32[7:0] ? content_249 : _GEN_2044; // @[Cat.scala 29:58]
  wire  _GEN_2046 = 8'hfa == _T_32[7:0] ? content_250 : _GEN_2045; // @[Cat.scala 29:58]
  wire  _GEN_2047 = 8'hfb == _T_32[7:0] ? content_251 : _GEN_2046; // @[Cat.scala 29:58]
  wire  _GEN_2048 = 8'hfc == _T_32[7:0] ? content_252 : _GEN_2047; // @[Cat.scala 29:58]
  wire  _GEN_2049 = 8'hfd == _T_32[7:0] ? content_253 : _GEN_2048; // @[Cat.scala 29:58]
  wire  _GEN_2050 = 8'hfe == _T_32[7:0] ? content_254 : _GEN_2049; // @[Cat.scala 29:58]
  wire  _GEN_2051 = 8'hff == _T_32[7:0] ? content_255 : _GEN_2050; // @[Cat.scala 29:58]
  wire  _GEN_2053 = 8'h1 == _T_42[7:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_2054 = 8'h2 == _T_42[7:0] ? content_2 : _GEN_2053; // @[Cat.scala 29:58]
  wire  _GEN_2055 = 8'h3 == _T_42[7:0] ? content_3 : _GEN_2054; // @[Cat.scala 29:58]
  wire  _GEN_2056 = 8'h4 == _T_42[7:0] ? content_4 : _GEN_2055; // @[Cat.scala 29:58]
  wire  _GEN_2057 = 8'h5 == _T_42[7:0] ? content_5 : _GEN_2056; // @[Cat.scala 29:58]
  wire  _GEN_2058 = 8'h6 == _T_42[7:0] ? content_6 : _GEN_2057; // @[Cat.scala 29:58]
  wire  _GEN_2059 = 8'h7 == _T_42[7:0] ? content_7 : _GEN_2058; // @[Cat.scala 29:58]
  wire  _GEN_2060 = 8'h8 == _T_42[7:0] ? content_8 : _GEN_2059; // @[Cat.scala 29:58]
  wire  _GEN_2061 = 8'h9 == _T_42[7:0] ? content_9 : _GEN_2060; // @[Cat.scala 29:58]
  wire  _GEN_2062 = 8'ha == _T_42[7:0] ? content_10 : _GEN_2061; // @[Cat.scala 29:58]
  wire  _GEN_2063 = 8'hb == _T_42[7:0] ? content_11 : _GEN_2062; // @[Cat.scala 29:58]
  wire  _GEN_2064 = 8'hc == _T_42[7:0] ? content_12 : _GEN_2063; // @[Cat.scala 29:58]
  wire  _GEN_2065 = 8'hd == _T_42[7:0] ? content_13 : _GEN_2064; // @[Cat.scala 29:58]
  wire  _GEN_2066 = 8'he == _T_42[7:0] ? content_14 : _GEN_2065; // @[Cat.scala 29:58]
  wire  _GEN_2067 = 8'hf == _T_42[7:0] ? content_15 : _GEN_2066; // @[Cat.scala 29:58]
  wire  _GEN_2068 = 8'h10 == _T_42[7:0] ? content_16 : _GEN_2067; // @[Cat.scala 29:58]
  wire  _GEN_2069 = 8'h11 == _T_42[7:0] ? content_17 : _GEN_2068; // @[Cat.scala 29:58]
  wire  _GEN_2070 = 8'h12 == _T_42[7:0] ? content_18 : _GEN_2069; // @[Cat.scala 29:58]
  wire  _GEN_2071 = 8'h13 == _T_42[7:0] ? content_19 : _GEN_2070; // @[Cat.scala 29:58]
  wire  _GEN_2072 = 8'h14 == _T_42[7:0] ? content_20 : _GEN_2071; // @[Cat.scala 29:58]
  wire  _GEN_2073 = 8'h15 == _T_42[7:0] ? content_21 : _GEN_2072; // @[Cat.scala 29:58]
  wire  _GEN_2074 = 8'h16 == _T_42[7:0] ? content_22 : _GEN_2073; // @[Cat.scala 29:58]
  wire  _GEN_2075 = 8'h17 == _T_42[7:0] ? content_23 : _GEN_2074; // @[Cat.scala 29:58]
  wire  _GEN_2076 = 8'h18 == _T_42[7:0] ? content_24 : _GEN_2075; // @[Cat.scala 29:58]
  wire  _GEN_2077 = 8'h19 == _T_42[7:0] ? content_25 : _GEN_2076; // @[Cat.scala 29:58]
  wire  _GEN_2078 = 8'h1a == _T_42[7:0] ? content_26 : _GEN_2077; // @[Cat.scala 29:58]
  wire  _GEN_2079 = 8'h1b == _T_42[7:0] ? content_27 : _GEN_2078; // @[Cat.scala 29:58]
  wire  _GEN_2080 = 8'h1c == _T_42[7:0] ? content_28 : _GEN_2079; // @[Cat.scala 29:58]
  wire  _GEN_2081 = 8'h1d == _T_42[7:0] ? content_29 : _GEN_2080; // @[Cat.scala 29:58]
  wire  _GEN_2082 = 8'h1e == _T_42[7:0] ? content_30 : _GEN_2081; // @[Cat.scala 29:58]
  wire  _GEN_2083 = 8'h1f == _T_42[7:0] ? content_31 : _GEN_2082; // @[Cat.scala 29:58]
  wire  _GEN_2084 = 8'h20 == _T_42[7:0] ? content_32 : _GEN_2083; // @[Cat.scala 29:58]
  wire  _GEN_2085 = 8'h21 == _T_42[7:0] ? content_33 : _GEN_2084; // @[Cat.scala 29:58]
  wire  _GEN_2086 = 8'h22 == _T_42[7:0] ? content_34 : _GEN_2085; // @[Cat.scala 29:58]
  wire  _GEN_2087 = 8'h23 == _T_42[7:0] ? content_35 : _GEN_2086; // @[Cat.scala 29:58]
  wire  _GEN_2088 = 8'h24 == _T_42[7:0] ? content_36 : _GEN_2087; // @[Cat.scala 29:58]
  wire  _GEN_2089 = 8'h25 == _T_42[7:0] ? content_37 : _GEN_2088; // @[Cat.scala 29:58]
  wire  _GEN_2090 = 8'h26 == _T_42[7:0] ? content_38 : _GEN_2089; // @[Cat.scala 29:58]
  wire  _GEN_2091 = 8'h27 == _T_42[7:0] ? content_39 : _GEN_2090; // @[Cat.scala 29:58]
  wire  _GEN_2092 = 8'h28 == _T_42[7:0] ? content_40 : _GEN_2091; // @[Cat.scala 29:58]
  wire  _GEN_2093 = 8'h29 == _T_42[7:0] ? content_41 : _GEN_2092; // @[Cat.scala 29:58]
  wire  _GEN_2094 = 8'h2a == _T_42[7:0] ? content_42 : _GEN_2093; // @[Cat.scala 29:58]
  wire  _GEN_2095 = 8'h2b == _T_42[7:0] ? content_43 : _GEN_2094; // @[Cat.scala 29:58]
  wire  _GEN_2096 = 8'h2c == _T_42[7:0] ? content_44 : _GEN_2095; // @[Cat.scala 29:58]
  wire  _GEN_2097 = 8'h2d == _T_42[7:0] ? content_45 : _GEN_2096; // @[Cat.scala 29:58]
  wire  _GEN_2098 = 8'h2e == _T_42[7:0] ? content_46 : _GEN_2097; // @[Cat.scala 29:58]
  wire  _GEN_2099 = 8'h2f == _T_42[7:0] ? content_47 : _GEN_2098; // @[Cat.scala 29:58]
  wire  _GEN_2100 = 8'h30 == _T_42[7:0] ? content_48 : _GEN_2099; // @[Cat.scala 29:58]
  wire  _GEN_2101 = 8'h31 == _T_42[7:0] ? content_49 : _GEN_2100; // @[Cat.scala 29:58]
  wire  _GEN_2102 = 8'h32 == _T_42[7:0] ? content_50 : _GEN_2101; // @[Cat.scala 29:58]
  wire  _GEN_2103 = 8'h33 == _T_42[7:0] ? content_51 : _GEN_2102; // @[Cat.scala 29:58]
  wire  _GEN_2104 = 8'h34 == _T_42[7:0] ? content_52 : _GEN_2103; // @[Cat.scala 29:58]
  wire  _GEN_2105 = 8'h35 == _T_42[7:0] ? content_53 : _GEN_2104; // @[Cat.scala 29:58]
  wire  _GEN_2106 = 8'h36 == _T_42[7:0] ? content_54 : _GEN_2105; // @[Cat.scala 29:58]
  wire  _GEN_2107 = 8'h37 == _T_42[7:0] ? content_55 : _GEN_2106; // @[Cat.scala 29:58]
  wire  _GEN_2108 = 8'h38 == _T_42[7:0] ? content_56 : _GEN_2107; // @[Cat.scala 29:58]
  wire  _GEN_2109 = 8'h39 == _T_42[7:0] ? content_57 : _GEN_2108; // @[Cat.scala 29:58]
  wire  _GEN_2110 = 8'h3a == _T_42[7:0] ? content_58 : _GEN_2109; // @[Cat.scala 29:58]
  wire  _GEN_2111 = 8'h3b == _T_42[7:0] ? content_59 : _GEN_2110; // @[Cat.scala 29:58]
  wire  _GEN_2112 = 8'h3c == _T_42[7:0] ? content_60 : _GEN_2111; // @[Cat.scala 29:58]
  wire  _GEN_2113 = 8'h3d == _T_42[7:0] ? content_61 : _GEN_2112; // @[Cat.scala 29:58]
  wire  _GEN_2114 = 8'h3e == _T_42[7:0] ? content_62 : _GEN_2113; // @[Cat.scala 29:58]
  wire  _GEN_2115 = 8'h3f == _T_42[7:0] ? content_63 : _GEN_2114; // @[Cat.scala 29:58]
  wire  _GEN_2116 = 8'h40 == _T_42[7:0] ? content_64 : _GEN_2115; // @[Cat.scala 29:58]
  wire  _GEN_2117 = 8'h41 == _T_42[7:0] ? content_65 : _GEN_2116; // @[Cat.scala 29:58]
  wire  _GEN_2118 = 8'h42 == _T_42[7:0] ? content_66 : _GEN_2117; // @[Cat.scala 29:58]
  wire  _GEN_2119 = 8'h43 == _T_42[7:0] ? content_67 : _GEN_2118; // @[Cat.scala 29:58]
  wire  _GEN_2120 = 8'h44 == _T_42[7:0] ? content_68 : _GEN_2119; // @[Cat.scala 29:58]
  wire  _GEN_2121 = 8'h45 == _T_42[7:0] ? content_69 : _GEN_2120; // @[Cat.scala 29:58]
  wire  _GEN_2122 = 8'h46 == _T_42[7:0] ? content_70 : _GEN_2121; // @[Cat.scala 29:58]
  wire  _GEN_2123 = 8'h47 == _T_42[7:0] ? content_71 : _GEN_2122; // @[Cat.scala 29:58]
  wire  _GEN_2124 = 8'h48 == _T_42[7:0] ? content_72 : _GEN_2123; // @[Cat.scala 29:58]
  wire  _GEN_2125 = 8'h49 == _T_42[7:0] ? content_73 : _GEN_2124; // @[Cat.scala 29:58]
  wire  _GEN_2126 = 8'h4a == _T_42[7:0] ? content_74 : _GEN_2125; // @[Cat.scala 29:58]
  wire  _GEN_2127 = 8'h4b == _T_42[7:0] ? content_75 : _GEN_2126; // @[Cat.scala 29:58]
  wire  _GEN_2128 = 8'h4c == _T_42[7:0] ? content_76 : _GEN_2127; // @[Cat.scala 29:58]
  wire  _GEN_2129 = 8'h4d == _T_42[7:0] ? content_77 : _GEN_2128; // @[Cat.scala 29:58]
  wire  _GEN_2130 = 8'h4e == _T_42[7:0] ? content_78 : _GEN_2129; // @[Cat.scala 29:58]
  wire  _GEN_2131 = 8'h4f == _T_42[7:0] ? content_79 : _GEN_2130; // @[Cat.scala 29:58]
  wire  _GEN_2132 = 8'h50 == _T_42[7:0] ? content_80 : _GEN_2131; // @[Cat.scala 29:58]
  wire  _GEN_2133 = 8'h51 == _T_42[7:0] ? content_81 : _GEN_2132; // @[Cat.scala 29:58]
  wire  _GEN_2134 = 8'h52 == _T_42[7:0] ? content_82 : _GEN_2133; // @[Cat.scala 29:58]
  wire  _GEN_2135 = 8'h53 == _T_42[7:0] ? content_83 : _GEN_2134; // @[Cat.scala 29:58]
  wire  _GEN_2136 = 8'h54 == _T_42[7:0] ? content_84 : _GEN_2135; // @[Cat.scala 29:58]
  wire  _GEN_2137 = 8'h55 == _T_42[7:0] ? content_85 : _GEN_2136; // @[Cat.scala 29:58]
  wire  _GEN_2138 = 8'h56 == _T_42[7:0] ? content_86 : _GEN_2137; // @[Cat.scala 29:58]
  wire  _GEN_2139 = 8'h57 == _T_42[7:0] ? content_87 : _GEN_2138; // @[Cat.scala 29:58]
  wire  _GEN_2140 = 8'h58 == _T_42[7:0] ? content_88 : _GEN_2139; // @[Cat.scala 29:58]
  wire  _GEN_2141 = 8'h59 == _T_42[7:0] ? content_89 : _GEN_2140; // @[Cat.scala 29:58]
  wire  _GEN_2142 = 8'h5a == _T_42[7:0] ? content_90 : _GEN_2141; // @[Cat.scala 29:58]
  wire  _GEN_2143 = 8'h5b == _T_42[7:0] ? content_91 : _GEN_2142; // @[Cat.scala 29:58]
  wire  _GEN_2144 = 8'h5c == _T_42[7:0] ? content_92 : _GEN_2143; // @[Cat.scala 29:58]
  wire  _GEN_2145 = 8'h5d == _T_42[7:0] ? content_93 : _GEN_2144; // @[Cat.scala 29:58]
  wire  _GEN_2146 = 8'h5e == _T_42[7:0] ? content_94 : _GEN_2145; // @[Cat.scala 29:58]
  wire  _GEN_2147 = 8'h5f == _T_42[7:0] ? content_95 : _GEN_2146; // @[Cat.scala 29:58]
  wire  _GEN_2148 = 8'h60 == _T_42[7:0] ? content_96 : _GEN_2147; // @[Cat.scala 29:58]
  wire  _GEN_2149 = 8'h61 == _T_42[7:0] ? content_97 : _GEN_2148; // @[Cat.scala 29:58]
  wire  _GEN_2150 = 8'h62 == _T_42[7:0] ? content_98 : _GEN_2149; // @[Cat.scala 29:58]
  wire  _GEN_2151 = 8'h63 == _T_42[7:0] ? content_99 : _GEN_2150; // @[Cat.scala 29:58]
  wire  _GEN_2152 = 8'h64 == _T_42[7:0] ? content_100 : _GEN_2151; // @[Cat.scala 29:58]
  wire  _GEN_2153 = 8'h65 == _T_42[7:0] ? content_101 : _GEN_2152; // @[Cat.scala 29:58]
  wire  _GEN_2154 = 8'h66 == _T_42[7:0] ? content_102 : _GEN_2153; // @[Cat.scala 29:58]
  wire  _GEN_2155 = 8'h67 == _T_42[7:0] ? content_103 : _GEN_2154; // @[Cat.scala 29:58]
  wire  _GEN_2156 = 8'h68 == _T_42[7:0] ? content_104 : _GEN_2155; // @[Cat.scala 29:58]
  wire  _GEN_2157 = 8'h69 == _T_42[7:0] ? content_105 : _GEN_2156; // @[Cat.scala 29:58]
  wire  _GEN_2158 = 8'h6a == _T_42[7:0] ? content_106 : _GEN_2157; // @[Cat.scala 29:58]
  wire  _GEN_2159 = 8'h6b == _T_42[7:0] ? content_107 : _GEN_2158; // @[Cat.scala 29:58]
  wire  _GEN_2160 = 8'h6c == _T_42[7:0] ? content_108 : _GEN_2159; // @[Cat.scala 29:58]
  wire  _GEN_2161 = 8'h6d == _T_42[7:0] ? content_109 : _GEN_2160; // @[Cat.scala 29:58]
  wire  _GEN_2162 = 8'h6e == _T_42[7:0] ? content_110 : _GEN_2161; // @[Cat.scala 29:58]
  wire  _GEN_2163 = 8'h6f == _T_42[7:0] ? content_111 : _GEN_2162; // @[Cat.scala 29:58]
  wire  _GEN_2164 = 8'h70 == _T_42[7:0] ? content_112 : _GEN_2163; // @[Cat.scala 29:58]
  wire  _GEN_2165 = 8'h71 == _T_42[7:0] ? content_113 : _GEN_2164; // @[Cat.scala 29:58]
  wire  _GEN_2166 = 8'h72 == _T_42[7:0] ? content_114 : _GEN_2165; // @[Cat.scala 29:58]
  wire  _GEN_2167 = 8'h73 == _T_42[7:0] ? content_115 : _GEN_2166; // @[Cat.scala 29:58]
  wire  _GEN_2168 = 8'h74 == _T_42[7:0] ? content_116 : _GEN_2167; // @[Cat.scala 29:58]
  wire  _GEN_2169 = 8'h75 == _T_42[7:0] ? content_117 : _GEN_2168; // @[Cat.scala 29:58]
  wire  _GEN_2170 = 8'h76 == _T_42[7:0] ? content_118 : _GEN_2169; // @[Cat.scala 29:58]
  wire  _GEN_2171 = 8'h77 == _T_42[7:0] ? content_119 : _GEN_2170; // @[Cat.scala 29:58]
  wire  _GEN_2172 = 8'h78 == _T_42[7:0] ? content_120 : _GEN_2171; // @[Cat.scala 29:58]
  wire  _GEN_2173 = 8'h79 == _T_42[7:0] ? content_121 : _GEN_2172; // @[Cat.scala 29:58]
  wire  _GEN_2174 = 8'h7a == _T_42[7:0] ? content_122 : _GEN_2173; // @[Cat.scala 29:58]
  wire  _GEN_2175 = 8'h7b == _T_42[7:0] ? content_123 : _GEN_2174; // @[Cat.scala 29:58]
  wire  _GEN_2176 = 8'h7c == _T_42[7:0] ? content_124 : _GEN_2175; // @[Cat.scala 29:58]
  wire  _GEN_2177 = 8'h7d == _T_42[7:0] ? content_125 : _GEN_2176; // @[Cat.scala 29:58]
  wire  _GEN_2178 = 8'h7e == _T_42[7:0] ? content_126 : _GEN_2177; // @[Cat.scala 29:58]
  wire  _GEN_2179 = 8'h7f == _T_42[7:0] ? content_127 : _GEN_2178; // @[Cat.scala 29:58]
  wire  _GEN_2180 = 8'h80 == _T_42[7:0] ? content_128 : _GEN_2179; // @[Cat.scala 29:58]
  wire  _GEN_2181 = 8'h81 == _T_42[7:0] ? content_129 : _GEN_2180; // @[Cat.scala 29:58]
  wire  _GEN_2182 = 8'h82 == _T_42[7:0] ? content_130 : _GEN_2181; // @[Cat.scala 29:58]
  wire  _GEN_2183 = 8'h83 == _T_42[7:0] ? content_131 : _GEN_2182; // @[Cat.scala 29:58]
  wire  _GEN_2184 = 8'h84 == _T_42[7:0] ? content_132 : _GEN_2183; // @[Cat.scala 29:58]
  wire  _GEN_2185 = 8'h85 == _T_42[7:0] ? content_133 : _GEN_2184; // @[Cat.scala 29:58]
  wire  _GEN_2186 = 8'h86 == _T_42[7:0] ? content_134 : _GEN_2185; // @[Cat.scala 29:58]
  wire  _GEN_2187 = 8'h87 == _T_42[7:0] ? content_135 : _GEN_2186; // @[Cat.scala 29:58]
  wire  _GEN_2188 = 8'h88 == _T_42[7:0] ? content_136 : _GEN_2187; // @[Cat.scala 29:58]
  wire  _GEN_2189 = 8'h89 == _T_42[7:0] ? content_137 : _GEN_2188; // @[Cat.scala 29:58]
  wire  _GEN_2190 = 8'h8a == _T_42[7:0] ? content_138 : _GEN_2189; // @[Cat.scala 29:58]
  wire  _GEN_2191 = 8'h8b == _T_42[7:0] ? content_139 : _GEN_2190; // @[Cat.scala 29:58]
  wire  _GEN_2192 = 8'h8c == _T_42[7:0] ? content_140 : _GEN_2191; // @[Cat.scala 29:58]
  wire  _GEN_2193 = 8'h8d == _T_42[7:0] ? content_141 : _GEN_2192; // @[Cat.scala 29:58]
  wire  _GEN_2194 = 8'h8e == _T_42[7:0] ? content_142 : _GEN_2193; // @[Cat.scala 29:58]
  wire  _GEN_2195 = 8'h8f == _T_42[7:0] ? content_143 : _GEN_2194; // @[Cat.scala 29:58]
  wire  _GEN_2196 = 8'h90 == _T_42[7:0] ? content_144 : _GEN_2195; // @[Cat.scala 29:58]
  wire  _GEN_2197 = 8'h91 == _T_42[7:0] ? content_145 : _GEN_2196; // @[Cat.scala 29:58]
  wire  _GEN_2198 = 8'h92 == _T_42[7:0] ? content_146 : _GEN_2197; // @[Cat.scala 29:58]
  wire  _GEN_2199 = 8'h93 == _T_42[7:0] ? content_147 : _GEN_2198; // @[Cat.scala 29:58]
  wire  _GEN_2200 = 8'h94 == _T_42[7:0] ? content_148 : _GEN_2199; // @[Cat.scala 29:58]
  wire  _GEN_2201 = 8'h95 == _T_42[7:0] ? content_149 : _GEN_2200; // @[Cat.scala 29:58]
  wire  _GEN_2202 = 8'h96 == _T_42[7:0] ? content_150 : _GEN_2201; // @[Cat.scala 29:58]
  wire  _GEN_2203 = 8'h97 == _T_42[7:0] ? content_151 : _GEN_2202; // @[Cat.scala 29:58]
  wire  _GEN_2204 = 8'h98 == _T_42[7:0] ? content_152 : _GEN_2203; // @[Cat.scala 29:58]
  wire  _GEN_2205 = 8'h99 == _T_42[7:0] ? content_153 : _GEN_2204; // @[Cat.scala 29:58]
  wire  _GEN_2206 = 8'h9a == _T_42[7:0] ? content_154 : _GEN_2205; // @[Cat.scala 29:58]
  wire  _GEN_2207 = 8'h9b == _T_42[7:0] ? content_155 : _GEN_2206; // @[Cat.scala 29:58]
  wire  _GEN_2208 = 8'h9c == _T_42[7:0] ? content_156 : _GEN_2207; // @[Cat.scala 29:58]
  wire  _GEN_2209 = 8'h9d == _T_42[7:0] ? content_157 : _GEN_2208; // @[Cat.scala 29:58]
  wire  _GEN_2210 = 8'h9e == _T_42[7:0] ? content_158 : _GEN_2209; // @[Cat.scala 29:58]
  wire  _GEN_2211 = 8'h9f == _T_42[7:0] ? content_159 : _GEN_2210; // @[Cat.scala 29:58]
  wire  _GEN_2212 = 8'ha0 == _T_42[7:0] ? content_160 : _GEN_2211; // @[Cat.scala 29:58]
  wire  _GEN_2213 = 8'ha1 == _T_42[7:0] ? content_161 : _GEN_2212; // @[Cat.scala 29:58]
  wire  _GEN_2214 = 8'ha2 == _T_42[7:0] ? content_162 : _GEN_2213; // @[Cat.scala 29:58]
  wire  _GEN_2215 = 8'ha3 == _T_42[7:0] ? content_163 : _GEN_2214; // @[Cat.scala 29:58]
  wire  _GEN_2216 = 8'ha4 == _T_42[7:0] ? content_164 : _GEN_2215; // @[Cat.scala 29:58]
  wire  _GEN_2217 = 8'ha5 == _T_42[7:0] ? content_165 : _GEN_2216; // @[Cat.scala 29:58]
  wire  _GEN_2218 = 8'ha6 == _T_42[7:0] ? content_166 : _GEN_2217; // @[Cat.scala 29:58]
  wire  _GEN_2219 = 8'ha7 == _T_42[7:0] ? content_167 : _GEN_2218; // @[Cat.scala 29:58]
  wire  _GEN_2220 = 8'ha8 == _T_42[7:0] ? content_168 : _GEN_2219; // @[Cat.scala 29:58]
  wire  _GEN_2221 = 8'ha9 == _T_42[7:0] ? content_169 : _GEN_2220; // @[Cat.scala 29:58]
  wire  _GEN_2222 = 8'haa == _T_42[7:0] ? content_170 : _GEN_2221; // @[Cat.scala 29:58]
  wire  _GEN_2223 = 8'hab == _T_42[7:0] ? content_171 : _GEN_2222; // @[Cat.scala 29:58]
  wire  _GEN_2224 = 8'hac == _T_42[7:0] ? content_172 : _GEN_2223; // @[Cat.scala 29:58]
  wire  _GEN_2225 = 8'had == _T_42[7:0] ? content_173 : _GEN_2224; // @[Cat.scala 29:58]
  wire  _GEN_2226 = 8'hae == _T_42[7:0] ? content_174 : _GEN_2225; // @[Cat.scala 29:58]
  wire  _GEN_2227 = 8'haf == _T_42[7:0] ? content_175 : _GEN_2226; // @[Cat.scala 29:58]
  wire  _GEN_2228 = 8'hb0 == _T_42[7:0] ? content_176 : _GEN_2227; // @[Cat.scala 29:58]
  wire  _GEN_2229 = 8'hb1 == _T_42[7:0] ? content_177 : _GEN_2228; // @[Cat.scala 29:58]
  wire  _GEN_2230 = 8'hb2 == _T_42[7:0] ? content_178 : _GEN_2229; // @[Cat.scala 29:58]
  wire  _GEN_2231 = 8'hb3 == _T_42[7:0] ? content_179 : _GEN_2230; // @[Cat.scala 29:58]
  wire  _GEN_2232 = 8'hb4 == _T_42[7:0] ? content_180 : _GEN_2231; // @[Cat.scala 29:58]
  wire  _GEN_2233 = 8'hb5 == _T_42[7:0] ? content_181 : _GEN_2232; // @[Cat.scala 29:58]
  wire  _GEN_2234 = 8'hb6 == _T_42[7:0] ? content_182 : _GEN_2233; // @[Cat.scala 29:58]
  wire  _GEN_2235 = 8'hb7 == _T_42[7:0] ? content_183 : _GEN_2234; // @[Cat.scala 29:58]
  wire  _GEN_2236 = 8'hb8 == _T_42[7:0] ? content_184 : _GEN_2235; // @[Cat.scala 29:58]
  wire  _GEN_2237 = 8'hb9 == _T_42[7:0] ? content_185 : _GEN_2236; // @[Cat.scala 29:58]
  wire  _GEN_2238 = 8'hba == _T_42[7:0] ? content_186 : _GEN_2237; // @[Cat.scala 29:58]
  wire  _GEN_2239 = 8'hbb == _T_42[7:0] ? content_187 : _GEN_2238; // @[Cat.scala 29:58]
  wire  _GEN_2240 = 8'hbc == _T_42[7:0] ? content_188 : _GEN_2239; // @[Cat.scala 29:58]
  wire  _GEN_2241 = 8'hbd == _T_42[7:0] ? content_189 : _GEN_2240; // @[Cat.scala 29:58]
  wire  _GEN_2242 = 8'hbe == _T_42[7:0] ? content_190 : _GEN_2241; // @[Cat.scala 29:58]
  wire  _GEN_2243 = 8'hbf == _T_42[7:0] ? content_191 : _GEN_2242; // @[Cat.scala 29:58]
  wire  _GEN_2244 = 8'hc0 == _T_42[7:0] ? content_192 : _GEN_2243; // @[Cat.scala 29:58]
  wire  _GEN_2245 = 8'hc1 == _T_42[7:0] ? content_193 : _GEN_2244; // @[Cat.scala 29:58]
  wire  _GEN_2246 = 8'hc2 == _T_42[7:0] ? content_194 : _GEN_2245; // @[Cat.scala 29:58]
  wire  _GEN_2247 = 8'hc3 == _T_42[7:0] ? content_195 : _GEN_2246; // @[Cat.scala 29:58]
  wire  _GEN_2248 = 8'hc4 == _T_42[7:0] ? content_196 : _GEN_2247; // @[Cat.scala 29:58]
  wire  _GEN_2249 = 8'hc5 == _T_42[7:0] ? content_197 : _GEN_2248; // @[Cat.scala 29:58]
  wire  _GEN_2250 = 8'hc6 == _T_42[7:0] ? content_198 : _GEN_2249; // @[Cat.scala 29:58]
  wire  _GEN_2251 = 8'hc7 == _T_42[7:0] ? content_199 : _GEN_2250; // @[Cat.scala 29:58]
  wire  _GEN_2252 = 8'hc8 == _T_42[7:0] ? content_200 : _GEN_2251; // @[Cat.scala 29:58]
  wire  _GEN_2253 = 8'hc9 == _T_42[7:0] ? content_201 : _GEN_2252; // @[Cat.scala 29:58]
  wire  _GEN_2254 = 8'hca == _T_42[7:0] ? content_202 : _GEN_2253; // @[Cat.scala 29:58]
  wire  _GEN_2255 = 8'hcb == _T_42[7:0] ? content_203 : _GEN_2254; // @[Cat.scala 29:58]
  wire  _GEN_2256 = 8'hcc == _T_42[7:0] ? content_204 : _GEN_2255; // @[Cat.scala 29:58]
  wire  _GEN_2257 = 8'hcd == _T_42[7:0] ? content_205 : _GEN_2256; // @[Cat.scala 29:58]
  wire  _GEN_2258 = 8'hce == _T_42[7:0] ? content_206 : _GEN_2257; // @[Cat.scala 29:58]
  wire  _GEN_2259 = 8'hcf == _T_42[7:0] ? content_207 : _GEN_2258; // @[Cat.scala 29:58]
  wire  _GEN_2260 = 8'hd0 == _T_42[7:0] ? content_208 : _GEN_2259; // @[Cat.scala 29:58]
  wire  _GEN_2261 = 8'hd1 == _T_42[7:0] ? content_209 : _GEN_2260; // @[Cat.scala 29:58]
  wire  _GEN_2262 = 8'hd2 == _T_42[7:0] ? content_210 : _GEN_2261; // @[Cat.scala 29:58]
  wire  _GEN_2263 = 8'hd3 == _T_42[7:0] ? content_211 : _GEN_2262; // @[Cat.scala 29:58]
  wire  _GEN_2264 = 8'hd4 == _T_42[7:0] ? content_212 : _GEN_2263; // @[Cat.scala 29:58]
  wire  _GEN_2265 = 8'hd5 == _T_42[7:0] ? content_213 : _GEN_2264; // @[Cat.scala 29:58]
  wire  _GEN_2266 = 8'hd6 == _T_42[7:0] ? content_214 : _GEN_2265; // @[Cat.scala 29:58]
  wire  _GEN_2267 = 8'hd7 == _T_42[7:0] ? content_215 : _GEN_2266; // @[Cat.scala 29:58]
  wire  _GEN_2268 = 8'hd8 == _T_42[7:0] ? content_216 : _GEN_2267; // @[Cat.scala 29:58]
  wire  _GEN_2269 = 8'hd9 == _T_42[7:0] ? content_217 : _GEN_2268; // @[Cat.scala 29:58]
  wire  _GEN_2270 = 8'hda == _T_42[7:0] ? content_218 : _GEN_2269; // @[Cat.scala 29:58]
  wire  _GEN_2271 = 8'hdb == _T_42[7:0] ? content_219 : _GEN_2270; // @[Cat.scala 29:58]
  wire  _GEN_2272 = 8'hdc == _T_42[7:0] ? content_220 : _GEN_2271; // @[Cat.scala 29:58]
  wire  _GEN_2273 = 8'hdd == _T_42[7:0] ? content_221 : _GEN_2272; // @[Cat.scala 29:58]
  wire  _GEN_2274 = 8'hde == _T_42[7:0] ? content_222 : _GEN_2273; // @[Cat.scala 29:58]
  wire  _GEN_2275 = 8'hdf == _T_42[7:0] ? content_223 : _GEN_2274; // @[Cat.scala 29:58]
  wire  _GEN_2276 = 8'he0 == _T_42[7:0] ? content_224 : _GEN_2275; // @[Cat.scala 29:58]
  wire  _GEN_2277 = 8'he1 == _T_42[7:0] ? content_225 : _GEN_2276; // @[Cat.scala 29:58]
  wire  _GEN_2278 = 8'he2 == _T_42[7:0] ? content_226 : _GEN_2277; // @[Cat.scala 29:58]
  wire  _GEN_2279 = 8'he3 == _T_42[7:0] ? content_227 : _GEN_2278; // @[Cat.scala 29:58]
  wire  _GEN_2280 = 8'he4 == _T_42[7:0] ? content_228 : _GEN_2279; // @[Cat.scala 29:58]
  wire  _GEN_2281 = 8'he5 == _T_42[7:0] ? content_229 : _GEN_2280; // @[Cat.scala 29:58]
  wire  _GEN_2282 = 8'he6 == _T_42[7:0] ? content_230 : _GEN_2281; // @[Cat.scala 29:58]
  wire  _GEN_2283 = 8'he7 == _T_42[7:0] ? content_231 : _GEN_2282; // @[Cat.scala 29:58]
  wire  _GEN_2284 = 8'he8 == _T_42[7:0] ? content_232 : _GEN_2283; // @[Cat.scala 29:58]
  wire  _GEN_2285 = 8'he9 == _T_42[7:0] ? content_233 : _GEN_2284; // @[Cat.scala 29:58]
  wire  _GEN_2286 = 8'hea == _T_42[7:0] ? content_234 : _GEN_2285; // @[Cat.scala 29:58]
  wire  _GEN_2287 = 8'heb == _T_42[7:0] ? content_235 : _GEN_2286; // @[Cat.scala 29:58]
  wire  _GEN_2288 = 8'hec == _T_42[7:0] ? content_236 : _GEN_2287; // @[Cat.scala 29:58]
  wire  _GEN_2289 = 8'hed == _T_42[7:0] ? content_237 : _GEN_2288; // @[Cat.scala 29:58]
  wire  _GEN_2290 = 8'hee == _T_42[7:0] ? content_238 : _GEN_2289; // @[Cat.scala 29:58]
  wire  _GEN_2291 = 8'hef == _T_42[7:0] ? content_239 : _GEN_2290; // @[Cat.scala 29:58]
  wire  _GEN_2292 = 8'hf0 == _T_42[7:0] ? content_240 : _GEN_2291; // @[Cat.scala 29:58]
  wire  _GEN_2293 = 8'hf1 == _T_42[7:0] ? content_241 : _GEN_2292; // @[Cat.scala 29:58]
  wire  _GEN_2294 = 8'hf2 == _T_42[7:0] ? content_242 : _GEN_2293; // @[Cat.scala 29:58]
  wire  _GEN_2295 = 8'hf3 == _T_42[7:0] ? content_243 : _GEN_2294; // @[Cat.scala 29:58]
  wire  _GEN_2296 = 8'hf4 == _T_42[7:0] ? content_244 : _GEN_2295; // @[Cat.scala 29:58]
  wire  _GEN_2297 = 8'hf5 == _T_42[7:0] ? content_245 : _GEN_2296; // @[Cat.scala 29:58]
  wire  _GEN_2298 = 8'hf6 == _T_42[7:0] ? content_246 : _GEN_2297; // @[Cat.scala 29:58]
  wire  _GEN_2299 = 8'hf7 == _T_42[7:0] ? content_247 : _GEN_2298; // @[Cat.scala 29:58]
  wire  _GEN_2300 = 8'hf8 == _T_42[7:0] ? content_248 : _GEN_2299; // @[Cat.scala 29:58]
  wire  _GEN_2301 = 8'hf9 == _T_42[7:0] ? content_249 : _GEN_2300; // @[Cat.scala 29:58]
  wire  _GEN_2302 = 8'hfa == _T_42[7:0] ? content_250 : _GEN_2301; // @[Cat.scala 29:58]
  wire  _GEN_2303 = 8'hfb == _T_42[7:0] ? content_251 : _GEN_2302; // @[Cat.scala 29:58]
  wire  _GEN_2304 = 8'hfc == _T_42[7:0] ? content_252 : _GEN_2303; // @[Cat.scala 29:58]
  wire  _GEN_2305 = 8'hfd == _T_42[7:0] ? content_253 : _GEN_2304; // @[Cat.scala 29:58]
  wire  _GEN_2306 = 8'hfe == _T_42[7:0] ? content_254 : _GEN_2305; // @[Cat.scala 29:58]
  wire  _GEN_2307 = 8'hff == _T_42[7:0] ? content_255 : _GEN_2306; // @[Cat.scala 29:58]
  wire  _GEN_2309 = 8'h1 == _T_39[7:0] ? content_1 : content_0; // @[Cat.scala 29:58]
  wire  _GEN_2310 = 8'h2 == _T_39[7:0] ? content_2 : _GEN_2309; // @[Cat.scala 29:58]
  wire  _GEN_2311 = 8'h3 == _T_39[7:0] ? content_3 : _GEN_2310; // @[Cat.scala 29:58]
  wire  _GEN_2312 = 8'h4 == _T_39[7:0] ? content_4 : _GEN_2311; // @[Cat.scala 29:58]
  wire  _GEN_2313 = 8'h5 == _T_39[7:0] ? content_5 : _GEN_2312; // @[Cat.scala 29:58]
  wire  _GEN_2314 = 8'h6 == _T_39[7:0] ? content_6 : _GEN_2313; // @[Cat.scala 29:58]
  wire  _GEN_2315 = 8'h7 == _T_39[7:0] ? content_7 : _GEN_2314; // @[Cat.scala 29:58]
  wire  _GEN_2316 = 8'h8 == _T_39[7:0] ? content_8 : _GEN_2315; // @[Cat.scala 29:58]
  wire  _GEN_2317 = 8'h9 == _T_39[7:0] ? content_9 : _GEN_2316; // @[Cat.scala 29:58]
  wire  _GEN_2318 = 8'ha == _T_39[7:0] ? content_10 : _GEN_2317; // @[Cat.scala 29:58]
  wire  _GEN_2319 = 8'hb == _T_39[7:0] ? content_11 : _GEN_2318; // @[Cat.scala 29:58]
  wire  _GEN_2320 = 8'hc == _T_39[7:0] ? content_12 : _GEN_2319; // @[Cat.scala 29:58]
  wire  _GEN_2321 = 8'hd == _T_39[7:0] ? content_13 : _GEN_2320; // @[Cat.scala 29:58]
  wire  _GEN_2322 = 8'he == _T_39[7:0] ? content_14 : _GEN_2321; // @[Cat.scala 29:58]
  wire  _GEN_2323 = 8'hf == _T_39[7:0] ? content_15 : _GEN_2322; // @[Cat.scala 29:58]
  wire  _GEN_2324 = 8'h10 == _T_39[7:0] ? content_16 : _GEN_2323; // @[Cat.scala 29:58]
  wire  _GEN_2325 = 8'h11 == _T_39[7:0] ? content_17 : _GEN_2324; // @[Cat.scala 29:58]
  wire  _GEN_2326 = 8'h12 == _T_39[7:0] ? content_18 : _GEN_2325; // @[Cat.scala 29:58]
  wire  _GEN_2327 = 8'h13 == _T_39[7:0] ? content_19 : _GEN_2326; // @[Cat.scala 29:58]
  wire  _GEN_2328 = 8'h14 == _T_39[7:0] ? content_20 : _GEN_2327; // @[Cat.scala 29:58]
  wire  _GEN_2329 = 8'h15 == _T_39[7:0] ? content_21 : _GEN_2328; // @[Cat.scala 29:58]
  wire  _GEN_2330 = 8'h16 == _T_39[7:0] ? content_22 : _GEN_2329; // @[Cat.scala 29:58]
  wire  _GEN_2331 = 8'h17 == _T_39[7:0] ? content_23 : _GEN_2330; // @[Cat.scala 29:58]
  wire  _GEN_2332 = 8'h18 == _T_39[7:0] ? content_24 : _GEN_2331; // @[Cat.scala 29:58]
  wire  _GEN_2333 = 8'h19 == _T_39[7:0] ? content_25 : _GEN_2332; // @[Cat.scala 29:58]
  wire  _GEN_2334 = 8'h1a == _T_39[7:0] ? content_26 : _GEN_2333; // @[Cat.scala 29:58]
  wire  _GEN_2335 = 8'h1b == _T_39[7:0] ? content_27 : _GEN_2334; // @[Cat.scala 29:58]
  wire  _GEN_2336 = 8'h1c == _T_39[7:0] ? content_28 : _GEN_2335; // @[Cat.scala 29:58]
  wire  _GEN_2337 = 8'h1d == _T_39[7:0] ? content_29 : _GEN_2336; // @[Cat.scala 29:58]
  wire  _GEN_2338 = 8'h1e == _T_39[7:0] ? content_30 : _GEN_2337; // @[Cat.scala 29:58]
  wire  _GEN_2339 = 8'h1f == _T_39[7:0] ? content_31 : _GEN_2338; // @[Cat.scala 29:58]
  wire  _GEN_2340 = 8'h20 == _T_39[7:0] ? content_32 : _GEN_2339; // @[Cat.scala 29:58]
  wire  _GEN_2341 = 8'h21 == _T_39[7:0] ? content_33 : _GEN_2340; // @[Cat.scala 29:58]
  wire  _GEN_2342 = 8'h22 == _T_39[7:0] ? content_34 : _GEN_2341; // @[Cat.scala 29:58]
  wire  _GEN_2343 = 8'h23 == _T_39[7:0] ? content_35 : _GEN_2342; // @[Cat.scala 29:58]
  wire  _GEN_2344 = 8'h24 == _T_39[7:0] ? content_36 : _GEN_2343; // @[Cat.scala 29:58]
  wire  _GEN_2345 = 8'h25 == _T_39[7:0] ? content_37 : _GEN_2344; // @[Cat.scala 29:58]
  wire  _GEN_2346 = 8'h26 == _T_39[7:0] ? content_38 : _GEN_2345; // @[Cat.scala 29:58]
  wire  _GEN_2347 = 8'h27 == _T_39[7:0] ? content_39 : _GEN_2346; // @[Cat.scala 29:58]
  wire  _GEN_2348 = 8'h28 == _T_39[7:0] ? content_40 : _GEN_2347; // @[Cat.scala 29:58]
  wire  _GEN_2349 = 8'h29 == _T_39[7:0] ? content_41 : _GEN_2348; // @[Cat.scala 29:58]
  wire  _GEN_2350 = 8'h2a == _T_39[7:0] ? content_42 : _GEN_2349; // @[Cat.scala 29:58]
  wire  _GEN_2351 = 8'h2b == _T_39[7:0] ? content_43 : _GEN_2350; // @[Cat.scala 29:58]
  wire  _GEN_2352 = 8'h2c == _T_39[7:0] ? content_44 : _GEN_2351; // @[Cat.scala 29:58]
  wire  _GEN_2353 = 8'h2d == _T_39[7:0] ? content_45 : _GEN_2352; // @[Cat.scala 29:58]
  wire  _GEN_2354 = 8'h2e == _T_39[7:0] ? content_46 : _GEN_2353; // @[Cat.scala 29:58]
  wire  _GEN_2355 = 8'h2f == _T_39[7:0] ? content_47 : _GEN_2354; // @[Cat.scala 29:58]
  wire  _GEN_2356 = 8'h30 == _T_39[7:0] ? content_48 : _GEN_2355; // @[Cat.scala 29:58]
  wire  _GEN_2357 = 8'h31 == _T_39[7:0] ? content_49 : _GEN_2356; // @[Cat.scala 29:58]
  wire  _GEN_2358 = 8'h32 == _T_39[7:0] ? content_50 : _GEN_2357; // @[Cat.scala 29:58]
  wire  _GEN_2359 = 8'h33 == _T_39[7:0] ? content_51 : _GEN_2358; // @[Cat.scala 29:58]
  wire  _GEN_2360 = 8'h34 == _T_39[7:0] ? content_52 : _GEN_2359; // @[Cat.scala 29:58]
  wire  _GEN_2361 = 8'h35 == _T_39[7:0] ? content_53 : _GEN_2360; // @[Cat.scala 29:58]
  wire  _GEN_2362 = 8'h36 == _T_39[7:0] ? content_54 : _GEN_2361; // @[Cat.scala 29:58]
  wire  _GEN_2363 = 8'h37 == _T_39[7:0] ? content_55 : _GEN_2362; // @[Cat.scala 29:58]
  wire  _GEN_2364 = 8'h38 == _T_39[7:0] ? content_56 : _GEN_2363; // @[Cat.scala 29:58]
  wire  _GEN_2365 = 8'h39 == _T_39[7:0] ? content_57 : _GEN_2364; // @[Cat.scala 29:58]
  wire  _GEN_2366 = 8'h3a == _T_39[7:0] ? content_58 : _GEN_2365; // @[Cat.scala 29:58]
  wire  _GEN_2367 = 8'h3b == _T_39[7:0] ? content_59 : _GEN_2366; // @[Cat.scala 29:58]
  wire  _GEN_2368 = 8'h3c == _T_39[7:0] ? content_60 : _GEN_2367; // @[Cat.scala 29:58]
  wire  _GEN_2369 = 8'h3d == _T_39[7:0] ? content_61 : _GEN_2368; // @[Cat.scala 29:58]
  wire  _GEN_2370 = 8'h3e == _T_39[7:0] ? content_62 : _GEN_2369; // @[Cat.scala 29:58]
  wire  _GEN_2371 = 8'h3f == _T_39[7:0] ? content_63 : _GEN_2370; // @[Cat.scala 29:58]
  wire  _GEN_2372 = 8'h40 == _T_39[7:0] ? content_64 : _GEN_2371; // @[Cat.scala 29:58]
  wire  _GEN_2373 = 8'h41 == _T_39[7:0] ? content_65 : _GEN_2372; // @[Cat.scala 29:58]
  wire  _GEN_2374 = 8'h42 == _T_39[7:0] ? content_66 : _GEN_2373; // @[Cat.scala 29:58]
  wire  _GEN_2375 = 8'h43 == _T_39[7:0] ? content_67 : _GEN_2374; // @[Cat.scala 29:58]
  wire  _GEN_2376 = 8'h44 == _T_39[7:0] ? content_68 : _GEN_2375; // @[Cat.scala 29:58]
  wire  _GEN_2377 = 8'h45 == _T_39[7:0] ? content_69 : _GEN_2376; // @[Cat.scala 29:58]
  wire  _GEN_2378 = 8'h46 == _T_39[7:0] ? content_70 : _GEN_2377; // @[Cat.scala 29:58]
  wire  _GEN_2379 = 8'h47 == _T_39[7:0] ? content_71 : _GEN_2378; // @[Cat.scala 29:58]
  wire  _GEN_2380 = 8'h48 == _T_39[7:0] ? content_72 : _GEN_2379; // @[Cat.scala 29:58]
  wire  _GEN_2381 = 8'h49 == _T_39[7:0] ? content_73 : _GEN_2380; // @[Cat.scala 29:58]
  wire  _GEN_2382 = 8'h4a == _T_39[7:0] ? content_74 : _GEN_2381; // @[Cat.scala 29:58]
  wire  _GEN_2383 = 8'h4b == _T_39[7:0] ? content_75 : _GEN_2382; // @[Cat.scala 29:58]
  wire  _GEN_2384 = 8'h4c == _T_39[7:0] ? content_76 : _GEN_2383; // @[Cat.scala 29:58]
  wire  _GEN_2385 = 8'h4d == _T_39[7:0] ? content_77 : _GEN_2384; // @[Cat.scala 29:58]
  wire  _GEN_2386 = 8'h4e == _T_39[7:0] ? content_78 : _GEN_2385; // @[Cat.scala 29:58]
  wire  _GEN_2387 = 8'h4f == _T_39[7:0] ? content_79 : _GEN_2386; // @[Cat.scala 29:58]
  wire  _GEN_2388 = 8'h50 == _T_39[7:0] ? content_80 : _GEN_2387; // @[Cat.scala 29:58]
  wire  _GEN_2389 = 8'h51 == _T_39[7:0] ? content_81 : _GEN_2388; // @[Cat.scala 29:58]
  wire  _GEN_2390 = 8'h52 == _T_39[7:0] ? content_82 : _GEN_2389; // @[Cat.scala 29:58]
  wire  _GEN_2391 = 8'h53 == _T_39[7:0] ? content_83 : _GEN_2390; // @[Cat.scala 29:58]
  wire  _GEN_2392 = 8'h54 == _T_39[7:0] ? content_84 : _GEN_2391; // @[Cat.scala 29:58]
  wire  _GEN_2393 = 8'h55 == _T_39[7:0] ? content_85 : _GEN_2392; // @[Cat.scala 29:58]
  wire  _GEN_2394 = 8'h56 == _T_39[7:0] ? content_86 : _GEN_2393; // @[Cat.scala 29:58]
  wire  _GEN_2395 = 8'h57 == _T_39[7:0] ? content_87 : _GEN_2394; // @[Cat.scala 29:58]
  wire  _GEN_2396 = 8'h58 == _T_39[7:0] ? content_88 : _GEN_2395; // @[Cat.scala 29:58]
  wire  _GEN_2397 = 8'h59 == _T_39[7:0] ? content_89 : _GEN_2396; // @[Cat.scala 29:58]
  wire  _GEN_2398 = 8'h5a == _T_39[7:0] ? content_90 : _GEN_2397; // @[Cat.scala 29:58]
  wire  _GEN_2399 = 8'h5b == _T_39[7:0] ? content_91 : _GEN_2398; // @[Cat.scala 29:58]
  wire  _GEN_2400 = 8'h5c == _T_39[7:0] ? content_92 : _GEN_2399; // @[Cat.scala 29:58]
  wire  _GEN_2401 = 8'h5d == _T_39[7:0] ? content_93 : _GEN_2400; // @[Cat.scala 29:58]
  wire  _GEN_2402 = 8'h5e == _T_39[7:0] ? content_94 : _GEN_2401; // @[Cat.scala 29:58]
  wire  _GEN_2403 = 8'h5f == _T_39[7:0] ? content_95 : _GEN_2402; // @[Cat.scala 29:58]
  wire  _GEN_2404 = 8'h60 == _T_39[7:0] ? content_96 : _GEN_2403; // @[Cat.scala 29:58]
  wire  _GEN_2405 = 8'h61 == _T_39[7:0] ? content_97 : _GEN_2404; // @[Cat.scala 29:58]
  wire  _GEN_2406 = 8'h62 == _T_39[7:0] ? content_98 : _GEN_2405; // @[Cat.scala 29:58]
  wire  _GEN_2407 = 8'h63 == _T_39[7:0] ? content_99 : _GEN_2406; // @[Cat.scala 29:58]
  wire  _GEN_2408 = 8'h64 == _T_39[7:0] ? content_100 : _GEN_2407; // @[Cat.scala 29:58]
  wire  _GEN_2409 = 8'h65 == _T_39[7:0] ? content_101 : _GEN_2408; // @[Cat.scala 29:58]
  wire  _GEN_2410 = 8'h66 == _T_39[7:0] ? content_102 : _GEN_2409; // @[Cat.scala 29:58]
  wire  _GEN_2411 = 8'h67 == _T_39[7:0] ? content_103 : _GEN_2410; // @[Cat.scala 29:58]
  wire  _GEN_2412 = 8'h68 == _T_39[7:0] ? content_104 : _GEN_2411; // @[Cat.scala 29:58]
  wire  _GEN_2413 = 8'h69 == _T_39[7:0] ? content_105 : _GEN_2412; // @[Cat.scala 29:58]
  wire  _GEN_2414 = 8'h6a == _T_39[7:0] ? content_106 : _GEN_2413; // @[Cat.scala 29:58]
  wire  _GEN_2415 = 8'h6b == _T_39[7:0] ? content_107 : _GEN_2414; // @[Cat.scala 29:58]
  wire  _GEN_2416 = 8'h6c == _T_39[7:0] ? content_108 : _GEN_2415; // @[Cat.scala 29:58]
  wire  _GEN_2417 = 8'h6d == _T_39[7:0] ? content_109 : _GEN_2416; // @[Cat.scala 29:58]
  wire  _GEN_2418 = 8'h6e == _T_39[7:0] ? content_110 : _GEN_2417; // @[Cat.scala 29:58]
  wire  _GEN_2419 = 8'h6f == _T_39[7:0] ? content_111 : _GEN_2418; // @[Cat.scala 29:58]
  wire  _GEN_2420 = 8'h70 == _T_39[7:0] ? content_112 : _GEN_2419; // @[Cat.scala 29:58]
  wire  _GEN_2421 = 8'h71 == _T_39[7:0] ? content_113 : _GEN_2420; // @[Cat.scala 29:58]
  wire  _GEN_2422 = 8'h72 == _T_39[7:0] ? content_114 : _GEN_2421; // @[Cat.scala 29:58]
  wire  _GEN_2423 = 8'h73 == _T_39[7:0] ? content_115 : _GEN_2422; // @[Cat.scala 29:58]
  wire  _GEN_2424 = 8'h74 == _T_39[7:0] ? content_116 : _GEN_2423; // @[Cat.scala 29:58]
  wire  _GEN_2425 = 8'h75 == _T_39[7:0] ? content_117 : _GEN_2424; // @[Cat.scala 29:58]
  wire  _GEN_2426 = 8'h76 == _T_39[7:0] ? content_118 : _GEN_2425; // @[Cat.scala 29:58]
  wire  _GEN_2427 = 8'h77 == _T_39[7:0] ? content_119 : _GEN_2426; // @[Cat.scala 29:58]
  wire  _GEN_2428 = 8'h78 == _T_39[7:0] ? content_120 : _GEN_2427; // @[Cat.scala 29:58]
  wire  _GEN_2429 = 8'h79 == _T_39[7:0] ? content_121 : _GEN_2428; // @[Cat.scala 29:58]
  wire  _GEN_2430 = 8'h7a == _T_39[7:0] ? content_122 : _GEN_2429; // @[Cat.scala 29:58]
  wire  _GEN_2431 = 8'h7b == _T_39[7:0] ? content_123 : _GEN_2430; // @[Cat.scala 29:58]
  wire  _GEN_2432 = 8'h7c == _T_39[7:0] ? content_124 : _GEN_2431; // @[Cat.scala 29:58]
  wire  _GEN_2433 = 8'h7d == _T_39[7:0] ? content_125 : _GEN_2432; // @[Cat.scala 29:58]
  wire  _GEN_2434 = 8'h7e == _T_39[7:0] ? content_126 : _GEN_2433; // @[Cat.scala 29:58]
  wire  _GEN_2435 = 8'h7f == _T_39[7:0] ? content_127 : _GEN_2434; // @[Cat.scala 29:58]
  wire  _GEN_2436 = 8'h80 == _T_39[7:0] ? content_128 : _GEN_2435; // @[Cat.scala 29:58]
  wire  _GEN_2437 = 8'h81 == _T_39[7:0] ? content_129 : _GEN_2436; // @[Cat.scala 29:58]
  wire  _GEN_2438 = 8'h82 == _T_39[7:0] ? content_130 : _GEN_2437; // @[Cat.scala 29:58]
  wire  _GEN_2439 = 8'h83 == _T_39[7:0] ? content_131 : _GEN_2438; // @[Cat.scala 29:58]
  wire  _GEN_2440 = 8'h84 == _T_39[7:0] ? content_132 : _GEN_2439; // @[Cat.scala 29:58]
  wire  _GEN_2441 = 8'h85 == _T_39[7:0] ? content_133 : _GEN_2440; // @[Cat.scala 29:58]
  wire  _GEN_2442 = 8'h86 == _T_39[7:0] ? content_134 : _GEN_2441; // @[Cat.scala 29:58]
  wire  _GEN_2443 = 8'h87 == _T_39[7:0] ? content_135 : _GEN_2442; // @[Cat.scala 29:58]
  wire  _GEN_2444 = 8'h88 == _T_39[7:0] ? content_136 : _GEN_2443; // @[Cat.scala 29:58]
  wire  _GEN_2445 = 8'h89 == _T_39[7:0] ? content_137 : _GEN_2444; // @[Cat.scala 29:58]
  wire  _GEN_2446 = 8'h8a == _T_39[7:0] ? content_138 : _GEN_2445; // @[Cat.scala 29:58]
  wire  _GEN_2447 = 8'h8b == _T_39[7:0] ? content_139 : _GEN_2446; // @[Cat.scala 29:58]
  wire  _GEN_2448 = 8'h8c == _T_39[7:0] ? content_140 : _GEN_2447; // @[Cat.scala 29:58]
  wire  _GEN_2449 = 8'h8d == _T_39[7:0] ? content_141 : _GEN_2448; // @[Cat.scala 29:58]
  wire  _GEN_2450 = 8'h8e == _T_39[7:0] ? content_142 : _GEN_2449; // @[Cat.scala 29:58]
  wire  _GEN_2451 = 8'h8f == _T_39[7:0] ? content_143 : _GEN_2450; // @[Cat.scala 29:58]
  wire  _GEN_2452 = 8'h90 == _T_39[7:0] ? content_144 : _GEN_2451; // @[Cat.scala 29:58]
  wire  _GEN_2453 = 8'h91 == _T_39[7:0] ? content_145 : _GEN_2452; // @[Cat.scala 29:58]
  wire  _GEN_2454 = 8'h92 == _T_39[7:0] ? content_146 : _GEN_2453; // @[Cat.scala 29:58]
  wire  _GEN_2455 = 8'h93 == _T_39[7:0] ? content_147 : _GEN_2454; // @[Cat.scala 29:58]
  wire  _GEN_2456 = 8'h94 == _T_39[7:0] ? content_148 : _GEN_2455; // @[Cat.scala 29:58]
  wire  _GEN_2457 = 8'h95 == _T_39[7:0] ? content_149 : _GEN_2456; // @[Cat.scala 29:58]
  wire  _GEN_2458 = 8'h96 == _T_39[7:0] ? content_150 : _GEN_2457; // @[Cat.scala 29:58]
  wire  _GEN_2459 = 8'h97 == _T_39[7:0] ? content_151 : _GEN_2458; // @[Cat.scala 29:58]
  wire  _GEN_2460 = 8'h98 == _T_39[7:0] ? content_152 : _GEN_2459; // @[Cat.scala 29:58]
  wire  _GEN_2461 = 8'h99 == _T_39[7:0] ? content_153 : _GEN_2460; // @[Cat.scala 29:58]
  wire  _GEN_2462 = 8'h9a == _T_39[7:0] ? content_154 : _GEN_2461; // @[Cat.scala 29:58]
  wire  _GEN_2463 = 8'h9b == _T_39[7:0] ? content_155 : _GEN_2462; // @[Cat.scala 29:58]
  wire  _GEN_2464 = 8'h9c == _T_39[7:0] ? content_156 : _GEN_2463; // @[Cat.scala 29:58]
  wire  _GEN_2465 = 8'h9d == _T_39[7:0] ? content_157 : _GEN_2464; // @[Cat.scala 29:58]
  wire  _GEN_2466 = 8'h9e == _T_39[7:0] ? content_158 : _GEN_2465; // @[Cat.scala 29:58]
  wire  _GEN_2467 = 8'h9f == _T_39[7:0] ? content_159 : _GEN_2466; // @[Cat.scala 29:58]
  wire  _GEN_2468 = 8'ha0 == _T_39[7:0] ? content_160 : _GEN_2467; // @[Cat.scala 29:58]
  wire  _GEN_2469 = 8'ha1 == _T_39[7:0] ? content_161 : _GEN_2468; // @[Cat.scala 29:58]
  wire  _GEN_2470 = 8'ha2 == _T_39[7:0] ? content_162 : _GEN_2469; // @[Cat.scala 29:58]
  wire  _GEN_2471 = 8'ha3 == _T_39[7:0] ? content_163 : _GEN_2470; // @[Cat.scala 29:58]
  wire  _GEN_2472 = 8'ha4 == _T_39[7:0] ? content_164 : _GEN_2471; // @[Cat.scala 29:58]
  wire  _GEN_2473 = 8'ha5 == _T_39[7:0] ? content_165 : _GEN_2472; // @[Cat.scala 29:58]
  wire  _GEN_2474 = 8'ha6 == _T_39[7:0] ? content_166 : _GEN_2473; // @[Cat.scala 29:58]
  wire  _GEN_2475 = 8'ha7 == _T_39[7:0] ? content_167 : _GEN_2474; // @[Cat.scala 29:58]
  wire  _GEN_2476 = 8'ha8 == _T_39[7:0] ? content_168 : _GEN_2475; // @[Cat.scala 29:58]
  wire  _GEN_2477 = 8'ha9 == _T_39[7:0] ? content_169 : _GEN_2476; // @[Cat.scala 29:58]
  wire  _GEN_2478 = 8'haa == _T_39[7:0] ? content_170 : _GEN_2477; // @[Cat.scala 29:58]
  wire  _GEN_2479 = 8'hab == _T_39[7:0] ? content_171 : _GEN_2478; // @[Cat.scala 29:58]
  wire  _GEN_2480 = 8'hac == _T_39[7:0] ? content_172 : _GEN_2479; // @[Cat.scala 29:58]
  wire  _GEN_2481 = 8'had == _T_39[7:0] ? content_173 : _GEN_2480; // @[Cat.scala 29:58]
  wire  _GEN_2482 = 8'hae == _T_39[7:0] ? content_174 : _GEN_2481; // @[Cat.scala 29:58]
  wire  _GEN_2483 = 8'haf == _T_39[7:0] ? content_175 : _GEN_2482; // @[Cat.scala 29:58]
  wire  _GEN_2484 = 8'hb0 == _T_39[7:0] ? content_176 : _GEN_2483; // @[Cat.scala 29:58]
  wire  _GEN_2485 = 8'hb1 == _T_39[7:0] ? content_177 : _GEN_2484; // @[Cat.scala 29:58]
  wire  _GEN_2486 = 8'hb2 == _T_39[7:0] ? content_178 : _GEN_2485; // @[Cat.scala 29:58]
  wire  _GEN_2487 = 8'hb3 == _T_39[7:0] ? content_179 : _GEN_2486; // @[Cat.scala 29:58]
  wire  _GEN_2488 = 8'hb4 == _T_39[7:0] ? content_180 : _GEN_2487; // @[Cat.scala 29:58]
  wire  _GEN_2489 = 8'hb5 == _T_39[7:0] ? content_181 : _GEN_2488; // @[Cat.scala 29:58]
  wire  _GEN_2490 = 8'hb6 == _T_39[7:0] ? content_182 : _GEN_2489; // @[Cat.scala 29:58]
  wire  _GEN_2491 = 8'hb7 == _T_39[7:0] ? content_183 : _GEN_2490; // @[Cat.scala 29:58]
  wire  _GEN_2492 = 8'hb8 == _T_39[7:0] ? content_184 : _GEN_2491; // @[Cat.scala 29:58]
  wire  _GEN_2493 = 8'hb9 == _T_39[7:0] ? content_185 : _GEN_2492; // @[Cat.scala 29:58]
  wire  _GEN_2494 = 8'hba == _T_39[7:0] ? content_186 : _GEN_2493; // @[Cat.scala 29:58]
  wire  _GEN_2495 = 8'hbb == _T_39[7:0] ? content_187 : _GEN_2494; // @[Cat.scala 29:58]
  wire  _GEN_2496 = 8'hbc == _T_39[7:0] ? content_188 : _GEN_2495; // @[Cat.scala 29:58]
  wire  _GEN_2497 = 8'hbd == _T_39[7:0] ? content_189 : _GEN_2496; // @[Cat.scala 29:58]
  wire  _GEN_2498 = 8'hbe == _T_39[7:0] ? content_190 : _GEN_2497; // @[Cat.scala 29:58]
  wire  _GEN_2499 = 8'hbf == _T_39[7:0] ? content_191 : _GEN_2498; // @[Cat.scala 29:58]
  wire  _GEN_2500 = 8'hc0 == _T_39[7:0] ? content_192 : _GEN_2499; // @[Cat.scala 29:58]
  wire  _GEN_2501 = 8'hc1 == _T_39[7:0] ? content_193 : _GEN_2500; // @[Cat.scala 29:58]
  wire  _GEN_2502 = 8'hc2 == _T_39[7:0] ? content_194 : _GEN_2501; // @[Cat.scala 29:58]
  wire  _GEN_2503 = 8'hc3 == _T_39[7:0] ? content_195 : _GEN_2502; // @[Cat.scala 29:58]
  wire  _GEN_2504 = 8'hc4 == _T_39[7:0] ? content_196 : _GEN_2503; // @[Cat.scala 29:58]
  wire  _GEN_2505 = 8'hc5 == _T_39[7:0] ? content_197 : _GEN_2504; // @[Cat.scala 29:58]
  wire  _GEN_2506 = 8'hc6 == _T_39[7:0] ? content_198 : _GEN_2505; // @[Cat.scala 29:58]
  wire  _GEN_2507 = 8'hc7 == _T_39[7:0] ? content_199 : _GEN_2506; // @[Cat.scala 29:58]
  wire  _GEN_2508 = 8'hc8 == _T_39[7:0] ? content_200 : _GEN_2507; // @[Cat.scala 29:58]
  wire  _GEN_2509 = 8'hc9 == _T_39[7:0] ? content_201 : _GEN_2508; // @[Cat.scala 29:58]
  wire  _GEN_2510 = 8'hca == _T_39[7:0] ? content_202 : _GEN_2509; // @[Cat.scala 29:58]
  wire  _GEN_2511 = 8'hcb == _T_39[7:0] ? content_203 : _GEN_2510; // @[Cat.scala 29:58]
  wire  _GEN_2512 = 8'hcc == _T_39[7:0] ? content_204 : _GEN_2511; // @[Cat.scala 29:58]
  wire  _GEN_2513 = 8'hcd == _T_39[7:0] ? content_205 : _GEN_2512; // @[Cat.scala 29:58]
  wire  _GEN_2514 = 8'hce == _T_39[7:0] ? content_206 : _GEN_2513; // @[Cat.scala 29:58]
  wire  _GEN_2515 = 8'hcf == _T_39[7:0] ? content_207 : _GEN_2514; // @[Cat.scala 29:58]
  wire  _GEN_2516 = 8'hd0 == _T_39[7:0] ? content_208 : _GEN_2515; // @[Cat.scala 29:58]
  wire  _GEN_2517 = 8'hd1 == _T_39[7:0] ? content_209 : _GEN_2516; // @[Cat.scala 29:58]
  wire  _GEN_2518 = 8'hd2 == _T_39[7:0] ? content_210 : _GEN_2517; // @[Cat.scala 29:58]
  wire  _GEN_2519 = 8'hd3 == _T_39[7:0] ? content_211 : _GEN_2518; // @[Cat.scala 29:58]
  wire  _GEN_2520 = 8'hd4 == _T_39[7:0] ? content_212 : _GEN_2519; // @[Cat.scala 29:58]
  wire  _GEN_2521 = 8'hd5 == _T_39[7:0] ? content_213 : _GEN_2520; // @[Cat.scala 29:58]
  wire  _GEN_2522 = 8'hd6 == _T_39[7:0] ? content_214 : _GEN_2521; // @[Cat.scala 29:58]
  wire  _GEN_2523 = 8'hd7 == _T_39[7:0] ? content_215 : _GEN_2522; // @[Cat.scala 29:58]
  wire  _GEN_2524 = 8'hd8 == _T_39[7:0] ? content_216 : _GEN_2523; // @[Cat.scala 29:58]
  wire  _GEN_2525 = 8'hd9 == _T_39[7:0] ? content_217 : _GEN_2524; // @[Cat.scala 29:58]
  wire  _GEN_2526 = 8'hda == _T_39[7:0] ? content_218 : _GEN_2525; // @[Cat.scala 29:58]
  wire  _GEN_2527 = 8'hdb == _T_39[7:0] ? content_219 : _GEN_2526; // @[Cat.scala 29:58]
  wire  _GEN_2528 = 8'hdc == _T_39[7:0] ? content_220 : _GEN_2527; // @[Cat.scala 29:58]
  wire  _GEN_2529 = 8'hdd == _T_39[7:0] ? content_221 : _GEN_2528; // @[Cat.scala 29:58]
  wire  _GEN_2530 = 8'hde == _T_39[7:0] ? content_222 : _GEN_2529; // @[Cat.scala 29:58]
  wire  _GEN_2531 = 8'hdf == _T_39[7:0] ? content_223 : _GEN_2530; // @[Cat.scala 29:58]
  wire  _GEN_2532 = 8'he0 == _T_39[7:0] ? content_224 : _GEN_2531; // @[Cat.scala 29:58]
  wire  _GEN_2533 = 8'he1 == _T_39[7:0] ? content_225 : _GEN_2532; // @[Cat.scala 29:58]
  wire  _GEN_2534 = 8'he2 == _T_39[7:0] ? content_226 : _GEN_2533; // @[Cat.scala 29:58]
  wire  _GEN_2535 = 8'he3 == _T_39[7:0] ? content_227 : _GEN_2534; // @[Cat.scala 29:58]
  wire  _GEN_2536 = 8'he4 == _T_39[7:0] ? content_228 : _GEN_2535; // @[Cat.scala 29:58]
  wire  _GEN_2537 = 8'he5 == _T_39[7:0] ? content_229 : _GEN_2536; // @[Cat.scala 29:58]
  wire  _GEN_2538 = 8'he6 == _T_39[7:0] ? content_230 : _GEN_2537; // @[Cat.scala 29:58]
  wire  _GEN_2539 = 8'he7 == _T_39[7:0] ? content_231 : _GEN_2538; // @[Cat.scala 29:58]
  wire  _GEN_2540 = 8'he8 == _T_39[7:0] ? content_232 : _GEN_2539; // @[Cat.scala 29:58]
  wire  _GEN_2541 = 8'he9 == _T_39[7:0] ? content_233 : _GEN_2540; // @[Cat.scala 29:58]
  wire  _GEN_2542 = 8'hea == _T_39[7:0] ? content_234 : _GEN_2541; // @[Cat.scala 29:58]
  wire  _GEN_2543 = 8'heb == _T_39[7:0] ? content_235 : _GEN_2542; // @[Cat.scala 29:58]
  wire  _GEN_2544 = 8'hec == _T_39[7:0] ? content_236 : _GEN_2543; // @[Cat.scala 29:58]
  wire  _GEN_2545 = 8'hed == _T_39[7:0] ? content_237 : _GEN_2544; // @[Cat.scala 29:58]
  wire  _GEN_2546 = 8'hee == _T_39[7:0] ? content_238 : _GEN_2545; // @[Cat.scala 29:58]
  wire  _GEN_2547 = 8'hef == _T_39[7:0] ? content_239 : _GEN_2546; // @[Cat.scala 29:58]
  wire  _GEN_2548 = 8'hf0 == _T_39[7:0] ? content_240 : _GEN_2547; // @[Cat.scala 29:58]
  wire  _GEN_2549 = 8'hf1 == _T_39[7:0] ? content_241 : _GEN_2548; // @[Cat.scala 29:58]
  wire  _GEN_2550 = 8'hf2 == _T_39[7:0] ? content_242 : _GEN_2549; // @[Cat.scala 29:58]
  wire  _GEN_2551 = 8'hf3 == _T_39[7:0] ? content_243 : _GEN_2550; // @[Cat.scala 29:58]
  wire  _GEN_2552 = 8'hf4 == _T_39[7:0] ? content_244 : _GEN_2551; // @[Cat.scala 29:58]
  wire  _GEN_2553 = 8'hf5 == _T_39[7:0] ? content_245 : _GEN_2552; // @[Cat.scala 29:58]
  wire  _GEN_2554 = 8'hf6 == _T_39[7:0] ? content_246 : _GEN_2553; // @[Cat.scala 29:58]
  wire  _GEN_2555 = 8'hf7 == _T_39[7:0] ? content_247 : _GEN_2554; // @[Cat.scala 29:58]
  wire  _GEN_2556 = 8'hf8 == _T_39[7:0] ? content_248 : _GEN_2555; // @[Cat.scala 29:58]
  wire  _GEN_2557 = 8'hf9 == _T_39[7:0] ? content_249 : _GEN_2556; // @[Cat.scala 29:58]
  wire  _GEN_2558 = 8'hfa == _T_39[7:0] ? content_250 : _GEN_2557; // @[Cat.scala 29:58]
  wire  _GEN_2559 = 8'hfb == _T_39[7:0] ? content_251 : _GEN_2558; // @[Cat.scala 29:58]
  wire  _GEN_2560 = 8'hfc == _T_39[7:0] ? content_252 : _GEN_2559; // @[Cat.scala 29:58]
  wire  _GEN_2561 = 8'hfd == _T_39[7:0] ? content_253 : _GEN_2560; // @[Cat.scala 29:58]
  wire  _GEN_2562 = 8'hfe == _T_39[7:0] ? content_254 : _GEN_2561; // @[Cat.scala 29:58]
  wire  _GEN_2563 = 8'hff == _T_39[7:0] ? content_255 : _GEN_2562; // @[Cat.scala 29:58]
  wire [3:0] _T_46 = {_GEN_2307,_GEN_2563,_GEN_1795,_GEN_2051}; // @[Cat.scala 29:58]
  assign io_port_0_read_out_0 = io_port_0_read_in_valid & _T_15[0]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_0_read_out_1 = io_port_0_read_in_valid & _T_15[1]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_0_read_out_2 = io_port_0_read_in_valid & _T_15[2]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_0_read_out_3 = io_port_0_read_in_valid & _T_15[3]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_1_read_out_0 = io_port_1_read_in_valid & _T_46[0]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_1_read_out_1 = io_port_1_read_in_valid & _T_46[1]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_1_read_out_2 = io_port_1_read_in_valid & _T_46[2]; // @[elements.scala 118:33 elements.scala 120:33]
  assign io_port_1_read_out_3 = io_port_1_read_in_valid & _T_46[3]; // @[elements.scala 118:33 elements.scala 120:33]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  content_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  content_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  content_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  content_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  content_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  content_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  content_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  content_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  content_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  content_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  content_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  content_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  content_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  content_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  content_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  content_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  content_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  content_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  content_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  content_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  content_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  content_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  content_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  content_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  content_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  content_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  content_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  content_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  content_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  content_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  content_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  content_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  content_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  content_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  content_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  content_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  content_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  content_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  content_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  content_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  content_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  content_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  content_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  content_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  content_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  content_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  content_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  content_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  content_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  content_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  content_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  content_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  content_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  content_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  content_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  content_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  content_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  content_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  content_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  content_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  content_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  content_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  content_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  content_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  content_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  content_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  content_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  content_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  content_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  content_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  content_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  content_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  content_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  content_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  content_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  content_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  content_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  content_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  content_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  content_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  content_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  content_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  content_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  content_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  content_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  content_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  content_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  content_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  content_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  content_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  content_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  content_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  content_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  content_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  content_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  content_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  content_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  content_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  content_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  content_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  content_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  content_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  content_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  content_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  content_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  content_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  content_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  content_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  content_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  content_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  content_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  content_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  content_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  content_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  content_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  content_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  content_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  content_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  content_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  content_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  content_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  content_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  content_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  content_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  content_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  content_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  content_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  content_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  content_128 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  content_129 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  content_130 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  content_131 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  content_132 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  content_133 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  content_134 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  content_135 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  content_136 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  content_137 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  content_138 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  content_139 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  content_140 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  content_141 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  content_142 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  content_143 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  content_144 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  content_145 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  content_146 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  content_147 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  content_148 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  content_149 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  content_150 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  content_151 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  content_152 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  content_153 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  content_154 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  content_155 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  content_156 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  content_157 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  content_158 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  content_159 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  content_160 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  content_161 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  content_162 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  content_163 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  content_164 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  content_165 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  content_166 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  content_167 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  content_168 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  content_169 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  content_170 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  content_171 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  content_172 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  content_173 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  content_174 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  content_175 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  content_176 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  content_177 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  content_178 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  content_179 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  content_180 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  content_181 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  content_182 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  content_183 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  content_184 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  content_185 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  content_186 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  content_187 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  content_188 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  content_189 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  content_190 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  content_191 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  content_192 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  content_193 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  content_194 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  content_195 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  content_196 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  content_197 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  content_198 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  content_199 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  content_200 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  content_201 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  content_202 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  content_203 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  content_204 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  content_205 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  content_206 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  content_207 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  content_208 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  content_209 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  content_210 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  content_211 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  content_212 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  content_213 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  content_214 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  content_215 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  content_216 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  content_217 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  content_218 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  content_219 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  content_220 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  content_221 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  content_222 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  content_223 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  content_224 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  content_225 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  content_226 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  content_227 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  content_228 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  content_229 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  content_230 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  content_231 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  content_232 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  content_233 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  content_234 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  content_235 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  content_236 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  content_237 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  content_238 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  content_239 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  content_240 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  content_241 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  content_242 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  content_243 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  content_244 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  content_245 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  content_246 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  content_247 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  content_248 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  content_249 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  content_250 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  content_251 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  content_252 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  content_253 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  content_254 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  content_255 = _RAND_255[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      content_0 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h0 == io_port_1_write_bits_addr[7:0]) begin
        content_0 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h0 == io_port_0_write_bits_addr[7:0]) begin
          content_0 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h0 == io_port_0_write_bits_addr[7:0]) begin
        content_0 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_1 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h1 == io_port_1_write_bits_addr[7:0]) begin
        content_1 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h1 == io_port_0_write_bits_addr[7:0]) begin
          content_1 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h1 == io_port_0_write_bits_addr[7:0]) begin
        content_1 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_2 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h2 == io_port_1_write_bits_addr[7:0]) begin
        content_2 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h2 == io_port_0_write_bits_addr[7:0]) begin
          content_2 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h2 == io_port_0_write_bits_addr[7:0]) begin
        content_2 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_3 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h3 == io_port_1_write_bits_addr[7:0]) begin
        content_3 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h3 == io_port_0_write_bits_addr[7:0]) begin
          content_3 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h3 == io_port_0_write_bits_addr[7:0]) begin
        content_3 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_4 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h4 == io_port_1_write_bits_addr[7:0]) begin
        content_4 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h4 == io_port_0_write_bits_addr[7:0]) begin
          content_4 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h4 == io_port_0_write_bits_addr[7:0]) begin
        content_4 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_5 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h5 == io_port_1_write_bits_addr[7:0]) begin
        content_5 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h5 == io_port_0_write_bits_addr[7:0]) begin
          content_5 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h5 == io_port_0_write_bits_addr[7:0]) begin
        content_5 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_6 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h6 == io_port_1_write_bits_addr[7:0]) begin
        content_6 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h6 == io_port_0_write_bits_addr[7:0]) begin
          content_6 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h6 == io_port_0_write_bits_addr[7:0]) begin
        content_6 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_7 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h7 == io_port_1_write_bits_addr[7:0]) begin
        content_7 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h7 == io_port_0_write_bits_addr[7:0]) begin
          content_7 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h7 == io_port_0_write_bits_addr[7:0]) begin
        content_7 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_8 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h8 == io_port_1_write_bits_addr[7:0]) begin
        content_8 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h8 == io_port_0_write_bits_addr[7:0]) begin
          content_8 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h8 == io_port_0_write_bits_addr[7:0]) begin
        content_8 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_9 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h9 == io_port_1_write_bits_addr[7:0]) begin
        content_9 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h9 == io_port_0_write_bits_addr[7:0]) begin
          content_9 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h9 == io_port_0_write_bits_addr[7:0]) begin
        content_9 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_10 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'ha == io_port_1_write_bits_addr[7:0]) begin
        content_10 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'ha == io_port_0_write_bits_addr[7:0]) begin
          content_10 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'ha == io_port_0_write_bits_addr[7:0]) begin
        content_10 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_11 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hb == io_port_1_write_bits_addr[7:0]) begin
        content_11 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hb == io_port_0_write_bits_addr[7:0]) begin
          content_11 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hb == io_port_0_write_bits_addr[7:0]) begin
        content_11 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_12 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hc == io_port_1_write_bits_addr[7:0]) begin
        content_12 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hc == io_port_0_write_bits_addr[7:0]) begin
          content_12 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hc == io_port_0_write_bits_addr[7:0]) begin
        content_12 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_13 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hd == io_port_1_write_bits_addr[7:0]) begin
        content_13 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hd == io_port_0_write_bits_addr[7:0]) begin
          content_13 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hd == io_port_0_write_bits_addr[7:0]) begin
        content_13 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_14 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'he == io_port_1_write_bits_addr[7:0]) begin
        content_14 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'he == io_port_0_write_bits_addr[7:0]) begin
          content_14 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'he == io_port_0_write_bits_addr[7:0]) begin
        content_14 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_15 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hf == io_port_1_write_bits_addr[7:0]) begin
        content_15 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hf == io_port_0_write_bits_addr[7:0]) begin
          content_15 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hf == io_port_0_write_bits_addr[7:0]) begin
        content_15 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_16 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h10 == io_port_1_write_bits_addr[7:0]) begin
        content_16 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h10 == io_port_0_write_bits_addr[7:0]) begin
          content_16 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h10 == io_port_0_write_bits_addr[7:0]) begin
        content_16 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_17 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h11 == io_port_1_write_bits_addr[7:0]) begin
        content_17 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h11 == io_port_0_write_bits_addr[7:0]) begin
          content_17 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h11 == io_port_0_write_bits_addr[7:0]) begin
        content_17 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_18 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h12 == io_port_1_write_bits_addr[7:0]) begin
        content_18 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h12 == io_port_0_write_bits_addr[7:0]) begin
          content_18 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h12 == io_port_0_write_bits_addr[7:0]) begin
        content_18 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_19 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h13 == io_port_1_write_bits_addr[7:0]) begin
        content_19 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h13 == io_port_0_write_bits_addr[7:0]) begin
          content_19 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h13 == io_port_0_write_bits_addr[7:0]) begin
        content_19 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_20 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h14 == io_port_1_write_bits_addr[7:0]) begin
        content_20 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h14 == io_port_0_write_bits_addr[7:0]) begin
          content_20 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h14 == io_port_0_write_bits_addr[7:0]) begin
        content_20 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_21 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h15 == io_port_1_write_bits_addr[7:0]) begin
        content_21 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h15 == io_port_0_write_bits_addr[7:0]) begin
          content_21 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h15 == io_port_0_write_bits_addr[7:0]) begin
        content_21 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_22 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h16 == io_port_1_write_bits_addr[7:0]) begin
        content_22 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h16 == io_port_0_write_bits_addr[7:0]) begin
          content_22 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h16 == io_port_0_write_bits_addr[7:0]) begin
        content_22 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_23 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h17 == io_port_1_write_bits_addr[7:0]) begin
        content_23 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h17 == io_port_0_write_bits_addr[7:0]) begin
          content_23 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h17 == io_port_0_write_bits_addr[7:0]) begin
        content_23 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_24 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h18 == io_port_1_write_bits_addr[7:0]) begin
        content_24 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h18 == io_port_0_write_bits_addr[7:0]) begin
          content_24 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h18 == io_port_0_write_bits_addr[7:0]) begin
        content_24 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_25 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h19 == io_port_1_write_bits_addr[7:0]) begin
        content_25 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h19 == io_port_0_write_bits_addr[7:0]) begin
          content_25 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h19 == io_port_0_write_bits_addr[7:0]) begin
        content_25 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_26 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h1a == io_port_1_write_bits_addr[7:0]) begin
        content_26 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h1a == io_port_0_write_bits_addr[7:0]) begin
          content_26 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h1a == io_port_0_write_bits_addr[7:0]) begin
        content_26 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_27 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h1b == io_port_1_write_bits_addr[7:0]) begin
        content_27 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h1b == io_port_0_write_bits_addr[7:0]) begin
          content_27 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h1b == io_port_0_write_bits_addr[7:0]) begin
        content_27 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_28 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h1c == io_port_1_write_bits_addr[7:0]) begin
        content_28 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h1c == io_port_0_write_bits_addr[7:0]) begin
          content_28 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h1c == io_port_0_write_bits_addr[7:0]) begin
        content_28 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_29 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h1d == io_port_1_write_bits_addr[7:0]) begin
        content_29 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h1d == io_port_0_write_bits_addr[7:0]) begin
          content_29 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h1d == io_port_0_write_bits_addr[7:0]) begin
        content_29 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_30 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h1e == io_port_1_write_bits_addr[7:0]) begin
        content_30 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h1e == io_port_0_write_bits_addr[7:0]) begin
          content_30 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h1e == io_port_0_write_bits_addr[7:0]) begin
        content_30 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_31 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h1f == io_port_1_write_bits_addr[7:0]) begin
        content_31 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h1f == io_port_0_write_bits_addr[7:0]) begin
          content_31 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h1f == io_port_0_write_bits_addr[7:0]) begin
        content_31 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_32 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h20 == io_port_1_write_bits_addr[7:0]) begin
        content_32 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h20 == io_port_0_write_bits_addr[7:0]) begin
          content_32 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h20 == io_port_0_write_bits_addr[7:0]) begin
        content_32 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_33 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h21 == io_port_1_write_bits_addr[7:0]) begin
        content_33 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h21 == io_port_0_write_bits_addr[7:0]) begin
          content_33 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h21 == io_port_0_write_bits_addr[7:0]) begin
        content_33 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_34 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h22 == io_port_1_write_bits_addr[7:0]) begin
        content_34 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h22 == io_port_0_write_bits_addr[7:0]) begin
          content_34 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h22 == io_port_0_write_bits_addr[7:0]) begin
        content_34 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_35 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h23 == io_port_1_write_bits_addr[7:0]) begin
        content_35 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h23 == io_port_0_write_bits_addr[7:0]) begin
          content_35 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h23 == io_port_0_write_bits_addr[7:0]) begin
        content_35 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_36 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h24 == io_port_1_write_bits_addr[7:0]) begin
        content_36 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h24 == io_port_0_write_bits_addr[7:0]) begin
          content_36 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h24 == io_port_0_write_bits_addr[7:0]) begin
        content_36 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_37 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h25 == io_port_1_write_bits_addr[7:0]) begin
        content_37 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h25 == io_port_0_write_bits_addr[7:0]) begin
          content_37 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h25 == io_port_0_write_bits_addr[7:0]) begin
        content_37 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_38 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h26 == io_port_1_write_bits_addr[7:0]) begin
        content_38 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h26 == io_port_0_write_bits_addr[7:0]) begin
          content_38 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h26 == io_port_0_write_bits_addr[7:0]) begin
        content_38 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_39 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h27 == io_port_1_write_bits_addr[7:0]) begin
        content_39 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h27 == io_port_0_write_bits_addr[7:0]) begin
          content_39 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h27 == io_port_0_write_bits_addr[7:0]) begin
        content_39 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_40 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h28 == io_port_1_write_bits_addr[7:0]) begin
        content_40 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h28 == io_port_0_write_bits_addr[7:0]) begin
          content_40 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h28 == io_port_0_write_bits_addr[7:0]) begin
        content_40 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_41 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h29 == io_port_1_write_bits_addr[7:0]) begin
        content_41 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h29 == io_port_0_write_bits_addr[7:0]) begin
          content_41 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h29 == io_port_0_write_bits_addr[7:0]) begin
        content_41 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_42 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h2a == io_port_1_write_bits_addr[7:0]) begin
        content_42 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h2a == io_port_0_write_bits_addr[7:0]) begin
          content_42 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h2a == io_port_0_write_bits_addr[7:0]) begin
        content_42 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_43 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h2b == io_port_1_write_bits_addr[7:0]) begin
        content_43 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h2b == io_port_0_write_bits_addr[7:0]) begin
          content_43 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h2b == io_port_0_write_bits_addr[7:0]) begin
        content_43 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_44 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h2c == io_port_1_write_bits_addr[7:0]) begin
        content_44 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h2c == io_port_0_write_bits_addr[7:0]) begin
          content_44 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h2c == io_port_0_write_bits_addr[7:0]) begin
        content_44 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_45 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h2d == io_port_1_write_bits_addr[7:0]) begin
        content_45 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h2d == io_port_0_write_bits_addr[7:0]) begin
          content_45 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h2d == io_port_0_write_bits_addr[7:0]) begin
        content_45 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_46 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h2e == io_port_1_write_bits_addr[7:0]) begin
        content_46 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h2e == io_port_0_write_bits_addr[7:0]) begin
          content_46 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h2e == io_port_0_write_bits_addr[7:0]) begin
        content_46 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_47 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h2f == io_port_1_write_bits_addr[7:0]) begin
        content_47 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h2f == io_port_0_write_bits_addr[7:0]) begin
          content_47 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h2f == io_port_0_write_bits_addr[7:0]) begin
        content_47 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_48 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h30 == io_port_1_write_bits_addr[7:0]) begin
        content_48 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h30 == io_port_0_write_bits_addr[7:0]) begin
          content_48 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h30 == io_port_0_write_bits_addr[7:0]) begin
        content_48 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_49 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h31 == io_port_1_write_bits_addr[7:0]) begin
        content_49 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h31 == io_port_0_write_bits_addr[7:0]) begin
          content_49 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h31 == io_port_0_write_bits_addr[7:0]) begin
        content_49 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_50 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h32 == io_port_1_write_bits_addr[7:0]) begin
        content_50 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h32 == io_port_0_write_bits_addr[7:0]) begin
          content_50 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h32 == io_port_0_write_bits_addr[7:0]) begin
        content_50 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_51 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h33 == io_port_1_write_bits_addr[7:0]) begin
        content_51 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h33 == io_port_0_write_bits_addr[7:0]) begin
          content_51 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h33 == io_port_0_write_bits_addr[7:0]) begin
        content_51 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_52 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h34 == io_port_1_write_bits_addr[7:0]) begin
        content_52 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h34 == io_port_0_write_bits_addr[7:0]) begin
          content_52 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h34 == io_port_0_write_bits_addr[7:0]) begin
        content_52 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_53 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h35 == io_port_1_write_bits_addr[7:0]) begin
        content_53 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h35 == io_port_0_write_bits_addr[7:0]) begin
          content_53 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h35 == io_port_0_write_bits_addr[7:0]) begin
        content_53 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_54 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h36 == io_port_1_write_bits_addr[7:0]) begin
        content_54 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h36 == io_port_0_write_bits_addr[7:0]) begin
          content_54 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h36 == io_port_0_write_bits_addr[7:0]) begin
        content_54 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_55 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h37 == io_port_1_write_bits_addr[7:0]) begin
        content_55 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h37 == io_port_0_write_bits_addr[7:0]) begin
          content_55 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h37 == io_port_0_write_bits_addr[7:0]) begin
        content_55 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_56 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h38 == io_port_1_write_bits_addr[7:0]) begin
        content_56 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h38 == io_port_0_write_bits_addr[7:0]) begin
          content_56 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h38 == io_port_0_write_bits_addr[7:0]) begin
        content_56 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_57 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h39 == io_port_1_write_bits_addr[7:0]) begin
        content_57 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h39 == io_port_0_write_bits_addr[7:0]) begin
          content_57 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h39 == io_port_0_write_bits_addr[7:0]) begin
        content_57 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_58 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h3a == io_port_1_write_bits_addr[7:0]) begin
        content_58 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h3a == io_port_0_write_bits_addr[7:0]) begin
          content_58 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h3a == io_port_0_write_bits_addr[7:0]) begin
        content_58 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_59 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h3b == io_port_1_write_bits_addr[7:0]) begin
        content_59 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h3b == io_port_0_write_bits_addr[7:0]) begin
          content_59 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h3b == io_port_0_write_bits_addr[7:0]) begin
        content_59 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_60 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h3c == io_port_1_write_bits_addr[7:0]) begin
        content_60 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h3c == io_port_0_write_bits_addr[7:0]) begin
          content_60 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h3c == io_port_0_write_bits_addr[7:0]) begin
        content_60 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_61 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h3d == io_port_1_write_bits_addr[7:0]) begin
        content_61 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h3d == io_port_0_write_bits_addr[7:0]) begin
          content_61 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h3d == io_port_0_write_bits_addr[7:0]) begin
        content_61 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_62 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h3e == io_port_1_write_bits_addr[7:0]) begin
        content_62 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h3e == io_port_0_write_bits_addr[7:0]) begin
          content_62 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h3e == io_port_0_write_bits_addr[7:0]) begin
        content_62 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_63 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h3f == io_port_1_write_bits_addr[7:0]) begin
        content_63 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h3f == io_port_0_write_bits_addr[7:0]) begin
          content_63 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h3f == io_port_0_write_bits_addr[7:0]) begin
        content_63 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_64 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h40 == io_port_1_write_bits_addr[7:0]) begin
        content_64 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h40 == io_port_0_write_bits_addr[7:0]) begin
          content_64 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h40 == io_port_0_write_bits_addr[7:0]) begin
        content_64 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_65 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h41 == io_port_1_write_bits_addr[7:0]) begin
        content_65 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h41 == io_port_0_write_bits_addr[7:0]) begin
          content_65 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h41 == io_port_0_write_bits_addr[7:0]) begin
        content_65 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_66 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h42 == io_port_1_write_bits_addr[7:0]) begin
        content_66 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h42 == io_port_0_write_bits_addr[7:0]) begin
          content_66 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h42 == io_port_0_write_bits_addr[7:0]) begin
        content_66 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_67 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h43 == io_port_1_write_bits_addr[7:0]) begin
        content_67 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h43 == io_port_0_write_bits_addr[7:0]) begin
          content_67 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h43 == io_port_0_write_bits_addr[7:0]) begin
        content_67 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_68 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h44 == io_port_1_write_bits_addr[7:0]) begin
        content_68 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h44 == io_port_0_write_bits_addr[7:0]) begin
          content_68 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h44 == io_port_0_write_bits_addr[7:0]) begin
        content_68 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_69 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h45 == io_port_1_write_bits_addr[7:0]) begin
        content_69 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h45 == io_port_0_write_bits_addr[7:0]) begin
          content_69 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h45 == io_port_0_write_bits_addr[7:0]) begin
        content_69 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_70 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h46 == io_port_1_write_bits_addr[7:0]) begin
        content_70 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h46 == io_port_0_write_bits_addr[7:0]) begin
          content_70 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h46 == io_port_0_write_bits_addr[7:0]) begin
        content_70 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_71 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h47 == io_port_1_write_bits_addr[7:0]) begin
        content_71 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h47 == io_port_0_write_bits_addr[7:0]) begin
          content_71 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h47 == io_port_0_write_bits_addr[7:0]) begin
        content_71 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_72 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h48 == io_port_1_write_bits_addr[7:0]) begin
        content_72 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h48 == io_port_0_write_bits_addr[7:0]) begin
          content_72 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h48 == io_port_0_write_bits_addr[7:0]) begin
        content_72 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_73 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h49 == io_port_1_write_bits_addr[7:0]) begin
        content_73 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h49 == io_port_0_write_bits_addr[7:0]) begin
          content_73 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h49 == io_port_0_write_bits_addr[7:0]) begin
        content_73 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_74 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h4a == io_port_1_write_bits_addr[7:0]) begin
        content_74 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h4a == io_port_0_write_bits_addr[7:0]) begin
          content_74 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h4a == io_port_0_write_bits_addr[7:0]) begin
        content_74 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_75 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h4b == io_port_1_write_bits_addr[7:0]) begin
        content_75 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h4b == io_port_0_write_bits_addr[7:0]) begin
          content_75 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h4b == io_port_0_write_bits_addr[7:0]) begin
        content_75 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_76 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h4c == io_port_1_write_bits_addr[7:0]) begin
        content_76 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h4c == io_port_0_write_bits_addr[7:0]) begin
          content_76 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h4c == io_port_0_write_bits_addr[7:0]) begin
        content_76 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_77 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h4d == io_port_1_write_bits_addr[7:0]) begin
        content_77 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h4d == io_port_0_write_bits_addr[7:0]) begin
          content_77 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h4d == io_port_0_write_bits_addr[7:0]) begin
        content_77 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_78 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h4e == io_port_1_write_bits_addr[7:0]) begin
        content_78 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h4e == io_port_0_write_bits_addr[7:0]) begin
          content_78 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h4e == io_port_0_write_bits_addr[7:0]) begin
        content_78 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_79 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h4f == io_port_1_write_bits_addr[7:0]) begin
        content_79 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h4f == io_port_0_write_bits_addr[7:0]) begin
          content_79 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h4f == io_port_0_write_bits_addr[7:0]) begin
        content_79 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_80 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h50 == io_port_1_write_bits_addr[7:0]) begin
        content_80 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h50 == io_port_0_write_bits_addr[7:0]) begin
          content_80 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h50 == io_port_0_write_bits_addr[7:0]) begin
        content_80 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_81 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h51 == io_port_1_write_bits_addr[7:0]) begin
        content_81 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h51 == io_port_0_write_bits_addr[7:0]) begin
          content_81 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h51 == io_port_0_write_bits_addr[7:0]) begin
        content_81 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_82 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h52 == io_port_1_write_bits_addr[7:0]) begin
        content_82 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h52 == io_port_0_write_bits_addr[7:0]) begin
          content_82 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h52 == io_port_0_write_bits_addr[7:0]) begin
        content_82 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_83 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h53 == io_port_1_write_bits_addr[7:0]) begin
        content_83 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h53 == io_port_0_write_bits_addr[7:0]) begin
          content_83 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h53 == io_port_0_write_bits_addr[7:0]) begin
        content_83 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_84 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h54 == io_port_1_write_bits_addr[7:0]) begin
        content_84 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h54 == io_port_0_write_bits_addr[7:0]) begin
          content_84 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h54 == io_port_0_write_bits_addr[7:0]) begin
        content_84 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_85 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h55 == io_port_1_write_bits_addr[7:0]) begin
        content_85 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h55 == io_port_0_write_bits_addr[7:0]) begin
          content_85 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h55 == io_port_0_write_bits_addr[7:0]) begin
        content_85 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_86 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h56 == io_port_1_write_bits_addr[7:0]) begin
        content_86 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h56 == io_port_0_write_bits_addr[7:0]) begin
          content_86 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h56 == io_port_0_write_bits_addr[7:0]) begin
        content_86 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_87 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h57 == io_port_1_write_bits_addr[7:0]) begin
        content_87 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h57 == io_port_0_write_bits_addr[7:0]) begin
          content_87 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h57 == io_port_0_write_bits_addr[7:0]) begin
        content_87 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_88 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h58 == io_port_1_write_bits_addr[7:0]) begin
        content_88 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h58 == io_port_0_write_bits_addr[7:0]) begin
          content_88 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h58 == io_port_0_write_bits_addr[7:0]) begin
        content_88 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_89 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h59 == io_port_1_write_bits_addr[7:0]) begin
        content_89 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h59 == io_port_0_write_bits_addr[7:0]) begin
          content_89 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h59 == io_port_0_write_bits_addr[7:0]) begin
        content_89 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_90 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h5a == io_port_1_write_bits_addr[7:0]) begin
        content_90 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h5a == io_port_0_write_bits_addr[7:0]) begin
          content_90 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h5a == io_port_0_write_bits_addr[7:0]) begin
        content_90 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_91 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h5b == io_port_1_write_bits_addr[7:0]) begin
        content_91 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h5b == io_port_0_write_bits_addr[7:0]) begin
          content_91 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h5b == io_port_0_write_bits_addr[7:0]) begin
        content_91 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_92 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h5c == io_port_1_write_bits_addr[7:0]) begin
        content_92 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h5c == io_port_0_write_bits_addr[7:0]) begin
          content_92 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h5c == io_port_0_write_bits_addr[7:0]) begin
        content_92 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_93 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h5d == io_port_1_write_bits_addr[7:0]) begin
        content_93 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h5d == io_port_0_write_bits_addr[7:0]) begin
          content_93 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h5d == io_port_0_write_bits_addr[7:0]) begin
        content_93 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_94 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h5e == io_port_1_write_bits_addr[7:0]) begin
        content_94 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h5e == io_port_0_write_bits_addr[7:0]) begin
          content_94 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h5e == io_port_0_write_bits_addr[7:0]) begin
        content_94 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_95 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h5f == io_port_1_write_bits_addr[7:0]) begin
        content_95 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h5f == io_port_0_write_bits_addr[7:0]) begin
          content_95 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h5f == io_port_0_write_bits_addr[7:0]) begin
        content_95 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_96 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h60 == io_port_1_write_bits_addr[7:0]) begin
        content_96 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h60 == io_port_0_write_bits_addr[7:0]) begin
          content_96 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h60 == io_port_0_write_bits_addr[7:0]) begin
        content_96 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_97 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h61 == io_port_1_write_bits_addr[7:0]) begin
        content_97 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h61 == io_port_0_write_bits_addr[7:0]) begin
          content_97 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h61 == io_port_0_write_bits_addr[7:0]) begin
        content_97 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_98 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h62 == io_port_1_write_bits_addr[7:0]) begin
        content_98 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h62 == io_port_0_write_bits_addr[7:0]) begin
          content_98 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h62 == io_port_0_write_bits_addr[7:0]) begin
        content_98 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_99 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h63 == io_port_1_write_bits_addr[7:0]) begin
        content_99 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h63 == io_port_0_write_bits_addr[7:0]) begin
          content_99 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h63 == io_port_0_write_bits_addr[7:0]) begin
        content_99 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_100 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h64 == io_port_1_write_bits_addr[7:0]) begin
        content_100 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h64 == io_port_0_write_bits_addr[7:0]) begin
          content_100 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h64 == io_port_0_write_bits_addr[7:0]) begin
        content_100 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_101 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h65 == io_port_1_write_bits_addr[7:0]) begin
        content_101 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h65 == io_port_0_write_bits_addr[7:0]) begin
          content_101 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h65 == io_port_0_write_bits_addr[7:0]) begin
        content_101 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_102 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h66 == io_port_1_write_bits_addr[7:0]) begin
        content_102 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h66 == io_port_0_write_bits_addr[7:0]) begin
          content_102 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h66 == io_port_0_write_bits_addr[7:0]) begin
        content_102 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_103 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h67 == io_port_1_write_bits_addr[7:0]) begin
        content_103 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h67 == io_port_0_write_bits_addr[7:0]) begin
          content_103 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h67 == io_port_0_write_bits_addr[7:0]) begin
        content_103 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_104 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h68 == io_port_1_write_bits_addr[7:0]) begin
        content_104 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h68 == io_port_0_write_bits_addr[7:0]) begin
          content_104 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h68 == io_port_0_write_bits_addr[7:0]) begin
        content_104 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_105 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h69 == io_port_1_write_bits_addr[7:0]) begin
        content_105 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h69 == io_port_0_write_bits_addr[7:0]) begin
          content_105 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h69 == io_port_0_write_bits_addr[7:0]) begin
        content_105 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_106 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h6a == io_port_1_write_bits_addr[7:0]) begin
        content_106 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h6a == io_port_0_write_bits_addr[7:0]) begin
          content_106 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h6a == io_port_0_write_bits_addr[7:0]) begin
        content_106 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_107 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h6b == io_port_1_write_bits_addr[7:0]) begin
        content_107 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h6b == io_port_0_write_bits_addr[7:0]) begin
          content_107 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h6b == io_port_0_write_bits_addr[7:0]) begin
        content_107 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_108 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h6c == io_port_1_write_bits_addr[7:0]) begin
        content_108 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h6c == io_port_0_write_bits_addr[7:0]) begin
          content_108 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h6c == io_port_0_write_bits_addr[7:0]) begin
        content_108 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_109 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h6d == io_port_1_write_bits_addr[7:0]) begin
        content_109 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h6d == io_port_0_write_bits_addr[7:0]) begin
          content_109 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h6d == io_port_0_write_bits_addr[7:0]) begin
        content_109 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_110 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h6e == io_port_1_write_bits_addr[7:0]) begin
        content_110 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h6e == io_port_0_write_bits_addr[7:0]) begin
          content_110 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h6e == io_port_0_write_bits_addr[7:0]) begin
        content_110 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_111 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h6f == io_port_1_write_bits_addr[7:0]) begin
        content_111 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h6f == io_port_0_write_bits_addr[7:0]) begin
          content_111 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h6f == io_port_0_write_bits_addr[7:0]) begin
        content_111 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_112 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h70 == io_port_1_write_bits_addr[7:0]) begin
        content_112 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h70 == io_port_0_write_bits_addr[7:0]) begin
          content_112 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h70 == io_port_0_write_bits_addr[7:0]) begin
        content_112 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_113 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h71 == io_port_1_write_bits_addr[7:0]) begin
        content_113 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h71 == io_port_0_write_bits_addr[7:0]) begin
          content_113 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h71 == io_port_0_write_bits_addr[7:0]) begin
        content_113 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_114 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h72 == io_port_1_write_bits_addr[7:0]) begin
        content_114 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h72 == io_port_0_write_bits_addr[7:0]) begin
          content_114 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h72 == io_port_0_write_bits_addr[7:0]) begin
        content_114 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_115 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h73 == io_port_1_write_bits_addr[7:0]) begin
        content_115 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h73 == io_port_0_write_bits_addr[7:0]) begin
          content_115 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h73 == io_port_0_write_bits_addr[7:0]) begin
        content_115 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_116 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h74 == io_port_1_write_bits_addr[7:0]) begin
        content_116 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h74 == io_port_0_write_bits_addr[7:0]) begin
          content_116 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h74 == io_port_0_write_bits_addr[7:0]) begin
        content_116 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_117 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h75 == io_port_1_write_bits_addr[7:0]) begin
        content_117 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h75 == io_port_0_write_bits_addr[7:0]) begin
          content_117 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h75 == io_port_0_write_bits_addr[7:0]) begin
        content_117 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_118 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h76 == io_port_1_write_bits_addr[7:0]) begin
        content_118 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h76 == io_port_0_write_bits_addr[7:0]) begin
          content_118 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h76 == io_port_0_write_bits_addr[7:0]) begin
        content_118 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_119 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h77 == io_port_1_write_bits_addr[7:0]) begin
        content_119 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h77 == io_port_0_write_bits_addr[7:0]) begin
          content_119 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h77 == io_port_0_write_bits_addr[7:0]) begin
        content_119 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_120 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h78 == io_port_1_write_bits_addr[7:0]) begin
        content_120 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h78 == io_port_0_write_bits_addr[7:0]) begin
          content_120 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h78 == io_port_0_write_bits_addr[7:0]) begin
        content_120 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_121 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h79 == io_port_1_write_bits_addr[7:0]) begin
        content_121 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h79 == io_port_0_write_bits_addr[7:0]) begin
          content_121 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h79 == io_port_0_write_bits_addr[7:0]) begin
        content_121 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_122 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h7a == io_port_1_write_bits_addr[7:0]) begin
        content_122 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h7a == io_port_0_write_bits_addr[7:0]) begin
          content_122 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h7a == io_port_0_write_bits_addr[7:0]) begin
        content_122 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_123 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h7b == io_port_1_write_bits_addr[7:0]) begin
        content_123 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h7b == io_port_0_write_bits_addr[7:0]) begin
          content_123 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h7b == io_port_0_write_bits_addr[7:0]) begin
        content_123 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_124 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h7c == io_port_1_write_bits_addr[7:0]) begin
        content_124 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h7c == io_port_0_write_bits_addr[7:0]) begin
          content_124 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h7c == io_port_0_write_bits_addr[7:0]) begin
        content_124 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_125 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h7d == io_port_1_write_bits_addr[7:0]) begin
        content_125 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h7d == io_port_0_write_bits_addr[7:0]) begin
          content_125 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h7d == io_port_0_write_bits_addr[7:0]) begin
        content_125 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_126 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h7e == io_port_1_write_bits_addr[7:0]) begin
        content_126 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h7e == io_port_0_write_bits_addr[7:0]) begin
          content_126 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h7e == io_port_0_write_bits_addr[7:0]) begin
        content_126 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_127 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h7f == io_port_1_write_bits_addr[7:0]) begin
        content_127 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h7f == io_port_0_write_bits_addr[7:0]) begin
          content_127 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h7f == io_port_0_write_bits_addr[7:0]) begin
        content_127 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_128 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h80 == io_port_1_write_bits_addr[7:0]) begin
        content_128 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h80 == io_port_0_write_bits_addr[7:0]) begin
          content_128 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h80 == io_port_0_write_bits_addr[7:0]) begin
        content_128 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_129 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h81 == io_port_1_write_bits_addr[7:0]) begin
        content_129 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h81 == io_port_0_write_bits_addr[7:0]) begin
          content_129 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h81 == io_port_0_write_bits_addr[7:0]) begin
        content_129 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_130 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h82 == io_port_1_write_bits_addr[7:0]) begin
        content_130 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h82 == io_port_0_write_bits_addr[7:0]) begin
          content_130 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h82 == io_port_0_write_bits_addr[7:0]) begin
        content_130 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_131 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h83 == io_port_1_write_bits_addr[7:0]) begin
        content_131 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h83 == io_port_0_write_bits_addr[7:0]) begin
          content_131 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h83 == io_port_0_write_bits_addr[7:0]) begin
        content_131 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_132 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h84 == io_port_1_write_bits_addr[7:0]) begin
        content_132 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h84 == io_port_0_write_bits_addr[7:0]) begin
          content_132 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h84 == io_port_0_write_bits_addr[7:0]) begin
        content_132 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_133 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h85 == io_port_1_write_bits_addr[7:0]) begin
        content_133 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h85 == io_port_0_write_bits_addr[7:0]) begin
          content_133 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h85 == io_port_0_write_bits_addr[7:0]) begin
        content_133 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_134 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h86 == io_port_1_write_bits_addr[7:0]) begin
        content_134 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h86 == io_port_0_write_bits_addr[7:0]) begin
          content_134 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h86 == io_port_0_write_bits_addr[7:0]) begin
        content_134 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_135 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h87 == io_port_1_write_bits_addr[7:0]) begin
        content_135 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h87 == io_port_0_write_bits_addr[7:0]) begin
          content_135 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h87 == io_port_0_write_bits_addr[7:0]) begin
        content_135 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_136 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h88 == io_port_1_write_bits_addr[7:0]) begin
        content_136 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h88 == io_port_0_write_bits_addr[7:0]) begin
          content_136 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h88 == io_port_0_write_bits_addr[7:0]) begin
        content_136 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_137 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h89 == io_port_1_write_bits_addr[7:0]) begin
        content_137 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h89 == io_port_0_write_bits_addr[7:0]) begin
          content_137 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h89 == io_port_0_write_bits_addr[7:0]) begin
        content_137 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_138 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h8a == io_port_1_write_bits_addr[7:0]) begin
        content_138 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h8a == io_port_0_write_bits_addr[7:0]) begin
          content_138 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h8a == io_port_0_write_bits_addr[7:0]) begin
        content_138 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_139 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h8b == io_port_1_write_bits_addr[7:0]) begin
        content_139 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h8b == io_port_0_write_bits_addr[7:0]) begin
          content_139 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h8b == io_port_0_write_bits_addr[7:0]) begin
        content_139 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_140 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h8c == io_port_1_write_bits_addr[7:0]) begin
        content_140 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h8c == io_port_0_write_bits_addr[7:0]) begin
          content_140 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h8c == io_port_0_write_bits_addr[7:0]) begin
        content_140 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_141 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h8d == io_port_1_write_bits_addr[7:0]) begin
        content_141 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h8d == io_port_0_write_bits_addr[7:0]) begin
          content_141 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h8d == io_port_0_write_bits_addr[7:0]) begin
        content_141 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_142 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h8e == io_port_1_write_bits_addr[7:0]) begin
        content_142 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h8e == io_port_0_write_bits_addr[7:0]) begin
          content_142 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h8e == io_port_0_write_bits_addr[7:0]) begin
        content_142 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_143 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h8f == io_port_1_write_bits_addr[7:0]) begin
        content_143 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h8f == io_port_0_write_bits_addr[7:0]) begin
          content_143 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h8f == io_port_0_write_bits_addr[7:0]) begin
        content_143 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_144 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h90 == io_port_1_write_bits_addr[7:0]) begin
        content_144 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h90 == io_port_0_write_bits_addr[7:0]) begin
          content_144 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h90 == io_port_0_write_bits_addr[7:0]) begin
        content_144 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_145 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h91 == io_port_1_write_bits_addr[7:0]) begin
        content_145 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h91 == io_port_0_write_bits_addr[7:0]) begin
          content_145 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h91 == io_port_0_write_bits_addr[7:0]) begin
        content_145 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_146 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h92 == io_port_1_write_bits_addr[7:0]) begin
        content_146 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h92 == io_port_0_write_bits_addr[7:0]) begin
          content_146 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h92 == io_port_0_write_bits_addr[7:0]) begin
        content_146 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_147 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h93 == io_port_1_write_bits_addr[7:0]) begin
        content_147 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h93 == io_port_0_write_bits_addr[7:0]) begin
          content_147 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h93 == io_port_0_write_bits_addr[7:0]) begin
        content_147 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_148 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h94 == io_port_1_write_bits_addr[7:0]) begin
        content_148 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h94 == io_port_0_write_bits_addr[7:0]) begin
          content_148 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h94 == io_port_0_write_bits_addr[7:0]) begin
        content_148 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_149 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h95 == io_port_1_write_bits_addr[7:0]) begin
        content_149 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h95 == io_port_0_write_bits_addr[7:0]) begin
          content_149 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h95 == io_port_0_write_bits_addr[7:0]) begin
        content_149 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_150 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h96 == io_port_1_write_bits_addr[7:0]) begin
        content_150 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h96 == io_port_0_write_bits_addr[7:0]) begin
          content_150 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h96 == io_port_0_write_bits_addr[7:0]) begin
        content_150 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_151 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h97 == io_port_1_write_bits_addr[7:0]) begin
        content_151 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h97 == io_port_0_write_bits_addr[7:0]) begin
          content_151 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h97 == io_port_0_write_bits_addr[7:0]) begin
        content_151 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_152 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h98 == io_port_1_write_bits_addr[7:0]) begin
        content_152 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h98 == io_port_0_write_bits_addr[7:0]) begin
          content_152 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h98 == io_port_0_write_bits_addr[7:0]) begin
        content_152 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_153 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h99 == io_port_1_write_bits_addr[7:0]) begin
        content_153 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h99 == io_port_0_write_bits_addr[7:0]) begin
          content_153 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h99 == io_port_0_write_bits_addr[7:0]) begin
        content_153 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_154 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h9a == io_port_1_write_bits_addr[7:0]) begin
        content_154 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h9a == io_port_0_write_bits_addr[7:0]) begin
          content_154 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h9a == io_port_0_write_bits_addr[7:0]) begin
        content_154 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_155 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h9b == io_port_1_write_bits_addr[7:0]) begin
        content_155 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h9b == io_port_0_write_bits_addr[7:0]) begin
          content_155 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h9b == io_port_0_write_bits_addr[7:0]) begin
        content_155 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_156 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h9c == io_port_1_write_bits_addr[7:0]) begin
        content_156 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h9c == io_port_0_write_bits_addr[7:0]) begin
          content_156 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h9c == io_port_0_write_bits_addr[7:0]) begin
        content_156 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_157 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h9d == io_port_1_write_bits_addr[7:0]) begin
        content_157 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h9d == io_port_0_write_bits_addr[7:0]) begin
          content_157 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h9d == io_port_0_write_bits_addr[7:0]) begin
        content_157 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_158 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h9e == io_port_1_write_bits_addr[7:0]) begin
        content_158 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h9e == io_port_0_write_bits_addr[7:0]) begin
          content_158 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h9e == io_port_0_write_bits_addr[7:0]) begin
        content_158 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_159 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'h9f == io_port_1_write_bits_addr[7:0]) begin
        content_159 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'h9f == io_port_0_write_bits_addr[7:0]) begin
          content_159 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'h9f == io_port_0_write_bits_addr[7:0]) begin
        content_159 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_160 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'ha0 == io_port_1_write_bits_addr[7:0]) begin
        content_160 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'ha0 == io_port_0_write_bits_addr[7:0]) begin
          content_160 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'ha0 == io_port_0_write_bits_addr[7:0]) begin
        content_160 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_161 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'ha1 == io_port_1_write_bits_addr[7:0]) begin
        content_161 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'ha1 == io_port_0_write_bits_addr[7:0]) begin
          content_161 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'ha1 == io_port_0_write_bits_addr[7:0]) begin
        content_161 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_162 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'ha2 == io_port_1_write_bits_addr[7:0]) begin
        content_162 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'ha2 == io_port_0_write_bits_addr[7:0]) begin
          content_162 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'ha2 == io_port_0_write_bits_addr[7:0]) begin
        content_162 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_163 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'ha3 == io_port_1_write_bits_addr[7:0]) begin
        content_163 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'ha3 == io_port_0_write_bits_addr[7:0]) begin
          content_163 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'ha3 == io_port_0_write_bits_addr[7:0]) begin
        content_163 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_164 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'ha4 == io_port_1_write_bits_addr[7:0]) begin
        content_164 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'ha4 == io_port_0_write_bits_addr[7:0]) begin
          content_164 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'ha4 == io_port_0_write_bits_addr[7:0]) begin
        content_164 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_165 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'ha5 == io_port_1_write_bits_addr[7:0]) begin
        content_165 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'ha5 == io_port_0_write_bits_addr[7:0]) begin
          content_165 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'ha5 == io_port_0_write_bits_addr[7:0]) begin
        content_165 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_166 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'ha6 == io_port_1_write_bits_addr[7:0]) begin
        content_166 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'ha6 == io_port_0_write_bits_addr[7:0]) begin
          content_166 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'ha6 == io_port_0_write_bits_addr[7:0]) begin
        content_166 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_167 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'ha7 == io_port_1_write_bits_addr[7:0]) begin
        content_167 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'ha7 == io_port_0_write_bits_addr[7:0]) begin
          content_167 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'ha7 == io_port_0_write_bits_addr[7:0]) begin
        content_167 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_168 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'ha8 == io_port_1_write_bits_addr[7:0]) begin
        content_168 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'ha8 == io_port_0_write_bits_addr[7:0]) begin
          content_168 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'ha8 == io_port_0_write_bits_addr[7:0]) begin
        content_168 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_169 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'ha9 == io_port_1_write_bits_addr[7:0]) begin
        content_169 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'ha9 == io_port_0_write_bits_addr[7:0]) begin
          content_169 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'ha9 == io_port_0_write_bits_addr[7:0]) begin
        content_169 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_170 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'haa == io_port_1_write_bits_addr[7:0]) begin
        content_170 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'haa == io_port_0_write_bits_addr[7:0]) begin
          content_170 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'haa == io_port_0_write_bits_addr[7:0]) begin
        content_170 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_171 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hab == io_port_1_write_bits_addr[7:0]) begin
        content_171 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hab == io_port_0_write_bits_addr[7:0]) begin
          content_171 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hab == io_port_0_write_bits_addr[7:0]) begin
        content_171 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_172 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hac == io_port_1_write_bits_addr[7:0]) begin
        content_172 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hac == io_port_0_write_bits_addr[7:0]) begin
          content_172 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hac == io_port_0_write_bits_addr[7:0]) begin
        content_172 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_173 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'had == io_port_1_write_bits_addr[7:0]) begin
        content_173 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'had == io_port_0_write_bits_addr[7:0]) begin
          content_173 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'had == io_port_0_write_bits_addr[7:0]) begin
        content_173 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_174 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hae == io_port_1_write_bits_addr[7:0]) begin
        content_174 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hae == io_port_0_write_bits_addr[7:0]) begin
          content_174 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hae == io_port_0_write_bits_addr[7:0]) begin
        content_174 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_175 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'haf == io_port_1_write_bits_addr[7:0]) begin
        content_175 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'haf == io_port_0_write_bits_addr[7:0]) begin
          content_175 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'haf == io_port_0_write_bits_addr[7:0]) begin
        content_175 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_176 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hb0 == io_port_1_write_bits_addr[7:0]) begin
        content_176 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hb0 == io_port_0_write_bits_addr[7:0]) begin
          content_176 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hb0 == io_port_0_write_bits_addr[7:0]) begin
        content_176 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_177 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hb1 == io_port_1_write_bits_addr[7:0]) begin
        content_177 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hb1 == io_port_0_write_bits_addr[7:0]) begin
          content_177 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hb1 == io_port_0_write_bits_addr[7:0]) begin
        content_177 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_178 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hb2 == io_port_1_write_bits_addr[7:0]) begin
        content_178 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hb2 == io_port_0_write_bits_addr[7:0]) begin
          content_178 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hb2 == io_port_0_write_bits_addr[7:0]) begin
        content_178 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_179 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hb3 == io_port_1_write_bits_addr[7:0]) begin
        content_179 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hb3 == io_port_0_write_bits_addr[7:0]) begin
          content_179 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hb3 == io_port_0_write_bits_addr[7:0]) begin
        content_179 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_180 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hb4 == io_port_1_write_bits_addr[7:0]) begin
        content_180 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hb4 == io_port_0_write_bits_addr[7:0]) begin
          content_180 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hb4 == io_port_0_write_bits_addr[7:0]) begin
        content_180 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_181 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hb5 == io_port_1_write_bits_addr[7:0]) begin
        content_181 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hb5 == io_port_0_write_bits_addr[7:0]) begin
          content_181 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hb5 == io_port_0_write_bits_addr[7:0]) begin
        content_181 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_182 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hb6 == io_port_1_write_bits_addr[7:0]) begin
        content_182 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hb6 == io_port_0_write_bits_addr[7:0]) begin
          content_182 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hb6 == io_port_0_write_bits_addr[7:0]) begin
        content_182 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_183 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hb7 == io_port_1_write_bits_addr[7:0]) begin
        content_183 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hb7 == io_port_0_write_bits_addr[7:0]) begin
          content_183 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hb7 == io_port_0_write_bits_addr[7:0]) begin
        content_183 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_184 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hb8 == io_port_1_write_bits_addr[7:0]) begin
        content_184 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hb8 == io_port_0_write_bits_addr[7:0]) begin
          content_184 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hb8 == io_port_0_write_bits_addr[7:0]) begin
        content_184 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_185 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hb9 == io_port_1_write_bits_addr[7:0]) begin
        content_185 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hb9 == io_port_0_write_bits_addr[7:0]) begin
          content_185 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hb9 == io_port_0_write_bits_addr[7:0]) begin
        content_185 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_186 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hba == io_port_1_write_bits_addr[7:0]) begin
        content_186 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hba == io_port_0_write_bits_addr[7:0]) begin
          content_186 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hba == io_port_0_write_bits_addr[7:0]) begin
        content_186 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_187 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hbb == io_port_1_write_bits_addr[7:0]) begin
        content_187 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hbb == io_port_0_write_bits_addr[7:0]) begin
          content_187 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hbb == io_port_0_write_bits_addr[7:0]) begin
        content_187 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_188 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hbc == io_port_1_write_bits_addr[7:0]) begin
        content_188 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hbc == io_port_0_write_bits_addr[7:0]) begin
          content_188 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hbc == io_port_0_write_bits_addr[7:0]) begin
        content_188 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_189 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hbd == io_port_1_write_bits_addr[7:0]) begin
        content_189 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hbd == io_port_0_write_bits_addr[7:0]) begin
          content_189 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hbd == io_port_0_write_bits_addr[7:0]) begin
        content_189 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_190 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hbe == io_port_1_write_bits_addr[7:0]) begin
        content_190 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hbe == io_port_0_write_bits_addr[7:0]) begin
          content_190 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hbe == io_port_0_write_bits_addr[7:0]) begin
        content_190 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_191 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hbf == io_port_1_write_bits_addr[7:0]) begin
        content_191 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hbf == io_port_0_write_bits_addr[7:0]) begin
          content_191 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hbf == io_port_0_write_bits_addr[7:0]) begin
        content_191 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_192 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hc0 == io_port_1_write_bits_addr[7:0]) begin
        content_192 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hc0 == io_port_0_write_bits_addr[7:0]) begin
          content_192 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hc0 == io_port_0_write_bits_addr[7:0]) begin
        content_192 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_193 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hc1 == io_port_1_write_bits_addr[7:0]) begin
        content_193 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hc1 == io_port_0_write_bits_addr[7:0]) begin
          content_193 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hc1 == io_port_0_write_bits_addr[7:0]) begin
        content_193 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_194 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hc2 == io_port_1_write_bits_addr[7:0]) begin
        content_194 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hc2 == io_port_0_write_bits_addr[7:0]) begin
          content_194 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hc2 == io_port_0_write_bits_addr[7:0]) begin
        content_194 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_195 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hc3 == io_port_1_write_bits_addr[7:0]) begin
        content_195 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hc3 == io_port_0_write_bits_addr[7:0]) begin
          content_195 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hc3 == io_port_0_write_bits_addr[7:0]) begin
        content_195 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_196 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hc4 == io_port_1_write_bits_addr[7:0]) begin
        content_196 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hc4 == io_port_0_write_bits_addr[7:0]) begin
          content_196 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hc4 == io_port_0_write_bits_addr[7:0]) begin
        content_196 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_197 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hc5 == io_port_1_write_bits_addr[7:0]) begin
        content_197 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hc5 == io_port_0_write_bits_addr[7:0]) begin
          content_197 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hc5 == io_port_0_write_bits_addr[7:0]) begin
        content_197 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_198 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hc6 == io_port_1_write_bits_addr[7:0]) begin
        content_198 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hc6 == io_port_0_write_bits_addr[7:0]) begin
          content_198 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hc6 == io_port_0_write_bits_addr[7:0]) begin
        content_198 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_199 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hc7 == io_port_1_write_bits_addr[7:0]) begin
        content_199 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hc7 == io_port_0_write_bits_addr[7:0]) begin
          content_199 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hc7 == io_port_0_write_bits_addr[7:0]) begin
        content_199 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_200 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hc8 == io_port_1_write_bits_addr[7:0]) begin
        content_200 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hc8 == io_port_0_write_bits_addr[7:0]) begin
          content_200 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hc8 == io_port_0_write_bits_addr[7:0]) begin
        content_200 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_201 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hc9 == io_port_1_write_bits_addr[7:0]) begin
        content_201 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hc9 == io_port_0_write_bits_addr[7:0]) begin
          content_201 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hc9 == io_port_0_write_bits_addr[7:0]) begin
        content_201 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_202 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hca == io_port_1_write_bits_addr[7:0]) begin
        content_202 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hca == io_port_0_write_bits_addr[7:0]) begin
          content_202 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hca == io_port_0_write_bits_addr[7:0]) begin
        content_202 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_203 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hcb == io_port_1_write_bits_addr[7:0]) begin
        content_203 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hcb == io_port_0_write_bits_addr[7:0]) begin
          content_203 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hcb == io_port_0_write_bits_addr[7:0]) begin
        content_203 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_204 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hcc == io_port_1_write_bits_addr[7:0]) begin
        content_204 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hcc == io_port_0_write_bits_addr[7:0]) begin
          content_204 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hcc == io_port_0_write_bits_addr[7:0]) begin
        content_204 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_205 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hcd == io_port_1_write_bits_addr[7:0]) begin
        content_205 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hcd == io_port_0_write_bits_addr[7:0]) begin
          content_205 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hcd == io_port_0_write_bits_addr[7:0]) begin
        content_205 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_206 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hce == io_port_1_write_bits_addr[7:0]) begin
        content_206 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hce == io_port_0_write_bits_addr[7:0]) begin
          content_206 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hce == io_port_0_write_bits_addr[7:0]) begin
        content_206 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_207 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hcf == io_port_1_write_bits_addr[7:0]) begin
        content_207 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hcf == io_port_0_write_bits_addr[7:0]) begin
          content_207 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hcf == io_port_0_write_bits_addr[7:0]) begin
        content_207 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_208 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hd0 == io_port_1_write_bits_addr[7:0]) begin
        content_208 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hd0 == io_port_0_write_bits_addr[7:0]) begin
          content_208 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hd0 == io_port_0_write_bits_addr[7:0]) begin
        content_208 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_209 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hd1 == io_port_1_write_bits_addr[7:0]) begin
        content_209 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hd1 == io_port_0_write_bits_addr[7:0]) begin
          content_209 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hd1 == io_port_0_write_bits_addr[7:0]) begin
        content_209 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_210 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hd2 == io_port_1_write_bits_addr[7:0]) begin
        content_210 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hd2 == io_port_0_write_bits_addr[7:0]) begin
          content_210 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hd2 == io_port_0_write_bits_addr[7:0]) begin
        content_210 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_211 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hd3 == io_port_1_write_bits_addr[7:0]) begin
        content_211 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hd3 == io_port_0_write_bits_addr[7:0]) begin
          content_211 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hd3 == io_port_0_write_bits_addr[7:0]) begin
        content_211 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_212 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hd4 == io_port_1_write_bits_addr[7:0]) begin
        content_212 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hd4 == io_port_0_write_bits_addr[7:0]) begin
          content_212 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hd4 == io_port_0_write_bits_addr[7:0]) begin
        content_212 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_213 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hd5 == io_port_1_write_bits_addr[7:0]) begin
        content_213 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hd5 == io_port_0_write_bits_addr[7:0]) begin
          content_213 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hd5 == io_port_0_write_bits_addr[7:0]) begin
        content_213 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_214 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hd6 == io_port_1_write_bits_addr[7:0]) begin
        content_214 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hd6 == io_port_0_write_bits_addr[7:0]) begin
          content_214 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hd6 == io_port_0_write_bits_addr[7:0]) begin
        content_214 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_215 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hd7 == io_port_1_write_bits_addr[7:0]) begin
        content_215 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hd7 == io_port_0_write_bits_addr[7:0]) begin
          content_215 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hd7 == io_port_0_write_bits_addr[7:0]) begin
        content_215 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_216 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hd8 == io_port_1_write_bits_addr[7:0]) begin
        content_216 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hd8 == io_port_0_write_bits_addr[7:0]) begin
          content_216 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hd8 == io_port_0_write_bits_addr[7:0]) begin
        content_216 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_217 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hd9 == io_port_1_write_bits_addr[7:0]) begin
        content_217 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hd9 == io_port_0_write_bits_addr[7:0]) begin
          content_217 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hd9 == io_port_0_write_bits_addr[7:0]) begin
        content_217 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_218 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hda == io_port_1_write_bits_addr[7:0]) begin
        content_218 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hda == io_port_0_write_bits_addr[7:0]) begin
          content_218 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hda == io_port_0_write_bits_addr[7:0]) begin
        content_218 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_219 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hdb == io_port_1_write_bits_addr[7:0]) begin
        content_219 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hdb == io_port_0_write_bits_addr[7:0]) begin
          content_219 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hdb == io_port_0_write_bits_addr[7:0]) begin
        content_219 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_220 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hdc == io_port_1_write_bits_addr[7:0]) begin
        content_220 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hdc == io_port_0_write_bits_addr[7:0]) begin
          content_220 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hdc == io_port_0_write_bits_addr[7:0]) begin
        content_220 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_221 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hdd == io_port_1_write_bits_addr[7:0]) begin
        content_221 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hdd == io_port_0_write_bits_addr[7:0]) begin
          content_221 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hdd == io_port_0_write_bits_addr[7:0]) begin
        content_221 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_222 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hde == io_port_1_write_bits_addr[7:0]) begin
        content_222 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hde == io_port_0_write_bits_addr[7:0]) begin
          content_222 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hde == io_port_0_write_bits_addr[7:0]) begin
        content_222 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_223 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hdf == io_port_1_write_bits_addr[7:0]) begin
        content_223 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hdf == io_port_0_write_bits_addr[7:0]) begin
          content_223 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hdf == io_port_0_write_bits_addr[7:0]) begin
        content_223 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_224 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'he0 == io_port_1_write_bits_addr[7:0]) begin
        content_224 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'he0 == io_port_0_write_bits_addr[7:0]) begin
          content_224 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'he0 == io_port_0_write_bits_addr[7:0]) begin
        content_224 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_225 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'he1 == io_port_1_write_bits_addr[7:0]) begin
        content_225 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'he1 == io_port_0_write_bits_addr[7:0]) begin
          content_225 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'he1 == io_port_0_write_bits_addr[7:0]) begin
        content_225 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_226 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'he2 == io_port_1_write_bits_addr[7:0]) begin
        content_226 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'he2 == io_port_0_write_bits_addr[7:0]) begin
          content_226 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'he2 == io_port_0_write_bits_addr[7:0]) begin
        content_226 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_227 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'he3 == io_port_1_write_bits_addr[7:0]) begin
        content_227 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'he3 == io_port_0_write_bits_addr[7:0]) begin
          content_227 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'he3 == io_port_0_write_bits_addr[7:0]) begin
        content_227 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_228 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'he4 == io_port_1_write_bits_addr[7:0]) begin
        content_228 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'he4 == io_port_0_write_bits_addr[7:0]) begin
          content_228 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'he4 == io_port_0_write_bits_addr[7:0]) begin
        content_228 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_229 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'he5 == io_port_1_write_bits_addr[7:0]) begin
        content_229 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'he5 == io_port_0_write_bits_addr[7:0]) begin
          content_229 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'he5 == io_port_0_write_bits_addr[7:0]) begin
        content_229 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_230 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'he6 == io_port_1_write_bits_addr[7:0]) begin
        content_230 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'he6 == io_port_0_write_bits_addr[7:0]) begin
          content_230 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'he6 == io_port_0_write_bits_addr[7:0]) begin
        content_230 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_231 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'he7 == io_port_1_write_bits_addr[7:0]) begin
        content_231 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'he7 == io_port_0_write_bits_addr[7:0]) begin
          content_231 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'he7 == io_port_0_write_bits_addr[7:0]) begin
        content_231 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_232 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'he8 == io_port_1_write_bits_addr[7:0]) begin
        content_232 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'he8 == io_port_0_write_bits_addr[7:0]) begin
          content_232 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'he8 == io_port_0_write_bits_addr[7:0]) begin
        content_232 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_233 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'he9 == io_port_1_write_bits_addr[7:0]) begin
        content_233 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'he9 == io_port_0_write_bits_addr[7:0]) begin
          content_233 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'he9 == io_port_0_write_bits_addr[7:0]) begin
        content_233 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_234 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hea == io_port_1_write_bits_addr[7:0]) begin
        content_234 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hea == io_port_0_write_bits_addr[7:0]) begin
          content_234 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hea == io_port_0_write_bits_addr[7:0]) begin
        content_234 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_235 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'heb == io_port_1_write_bits_addr[7:0]) begin
        content_235 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'heb == io_port_0_write_bits_addr[7:0]) begin
          content_235 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'heb == io_port_0_write_bits_addr[7:0]) begin
        content_235 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_236 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hec == io_port_1_write_bits_addr[7:0]) begin
        content_236 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hec == io_port_0_write_bits_addr[7:0]) begin
          content_236 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hec == io_port_0_write_bits_addr[7:0]) begin
        content_236 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_237 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hed == io_port_1_write_bits_addr[7:0]) begin
        content_237 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hed == io_port_0_write_bits_addr[7:0]) begin
          content_237 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hed == io_port_0_write_bits_addr[7:0]) begin
        content_237 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_238 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hee == io_port_1_write_bits_addr[7:0]) begin
        content_238 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hee == io_port_0_write_bits_addr[7:0]) begin
          content_238 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hee == io_port_0_write_bits_addr[7:0]) begin
        content_238 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_239 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hef == io_port_1_write_bits_addr[7:0]) begin
        content_239 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hef == io_port_0_write_bits_addr[7:0]) begin
          content_239 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hef == io_port_0_write_bits_addr[7:0]) begin
        content_239 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_240 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hf0 == io_port_1_write_bits_addr[7:0]) begin
        content_240 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hf0 == io_port_0_write_bits_addr[7:0]) begin
          content_240 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hf0 == io_port_0_write_bits_addr[7:0]) begin
        content_240 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_241 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hf1 == io_port_1_write_bits_addr[7:0]) begin
        content_241 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hf1 == io_port_0_write_bits_addr[7:0]) begin
          content_241 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hf1 == io_port_0_write_bits_addr[7:0]) begin
        content_241 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_242 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hf2 == io_port_1_write_bits_addr[7:0]) begin
        content_242 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hf2 == io_port_0_write_bits_addr[7:0]) begin
          content_242 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hf2 == io_port_0_write_bits_addr[7:0]) begin
        content_242 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_243 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hf3 == io_port_1_write_bits_addr[7:0]) begin
        content_243 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hf3 == io_port_0_write_bits_addr[7:0]) begin
          content_243 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hf3 == io_port_0_write_bits_addr[7:0]) begin
        content_243 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_244 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hf4 == io_port_1_write_bits_addr[7:0]) begin
        content_244 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hf4 == io_port_0_write_bits_addr[7:0]) begin
          content_244 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hf4 == io_port_0_write_bits_addr[7:0]) begin
        content_244 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_245 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hf5 == io_port_1_write_bits_addr[7:0]) begin
        content_245 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hf5 == io_port_0_write_bits_addr[7:0]) begin
          content_245 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hf5 == io_port_0_write_bits_addr[7:0]) begin
        content_245 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_246 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hf6 == io_port_1_write_bits_addr[7:0]) begin
        content_246 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hf6 == io_port_0_write_bits_addr[7:0]) begin
          content_246 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hf6 == io_port_0_write_bits_addr[7:0]) begin
        content_246 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_247 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hf7 == io_port_1_write_bits_addr[7:0]) begin
        content_247 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hf7 == io_port_0_write_bits_addr[7:0]) begin
          content_247 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hf7 == io_port_0_write_bits_addr[7:0]) begin
        content_247 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_248 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hf8 == io_port_1_write_bits_addr[7:0]) begin
        content_248 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hf8 == io_port_0_write_bits_addr[7:0]) begin
          content_248 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hf8 == io_port_0_write_bits_addr[7:0]) begin
        content_248 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_249 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hf9 == io_port_1_write_bits_addr[7:0]) begin
        content_249 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hf9 == io_port_0_write_bits_addr[7:0]) begin
          content_249 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hf9 == io_port_0_write_bits_addr[7:0]) begin
        content_249 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_250 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hfa == io_port_1_write_bits_addr[7:0]) begin
        content_250 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hfa == io_port_0_write_bits_addr[7:0]) begin
          content_250 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hfa == io_port_0_write_bits_addr[7:0]) begin
        content_250 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_251 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hfb == io_port_1_write_bits_addr[7:0]) begin
        content_251 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hfb == io_port_0_write_bits_addr[7:0]) begin
          content_251 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hfb == io_port_0_write_bits_addr[7:0]) begin
        content_251 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_252 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hfc == io_port_1_write_bits_addr[7:0]) begin
        content_252 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hfc == io_port_0_write_bits_addr[7:0]) begin
          content_252 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hfc == io_port_0_write_bits_addr[7:0]) begin
        content_252 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_253 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hfd == io_port_1_write_bits_addr[7:0]) begin
        content_253 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hfd == io_port_0_write_bits_addr[7:0]) begin
          content_253 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hfd == io_port_0_write_bits_addr[7:0]) begin
        content_253 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_254 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hfe == io_port_1_write_bits_addr[7:0]) begin
        content_254 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hfe == io_port_0_write_bits_addr[7:0]) begin
          content_254 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hfe == io_port_0_write_bits_addr[7:0]) begin
        content_254 <= io_port_0_write_bits_value;
      end
    end
    if (reset) begin
      content_255 <= 1'h0;
    end else if (io_port_1_write_valid) begin
      if (8'hff == io_port_1_write_bits_addr[7:0]) begin
        content_255 <= io_port_1_write_bits_value;
      end else if (io_port_0_write_valid) begin
        if (8'hff == io_port_0_write_bits_addr[7:0]) begin
          content_255 <= io_port_0_write_bits_value;
        end
      end
    end else if (io_port_0_write_valid) begin
      if (8'hff == io_port_0_write_bits_addr[7:0]) begin
        content_255 <= io_port_0_write_bits_value;
      end
    end
  end
endmodule
module Arbiter_2(
  input         io_in_0_valid,
  input  [3:0]  io_in_0_bits_bank,
  input  [5:0]  io_in_0_bits_address,
  input  [22:0] io_in_0_bits_inputValue_0_tag,
  input  [22:0] io_in_0_bits_inputValue_1_tag,
  input  [22:0] io_in_0_bits_inputValue_2_tag,
  input  [22:0] io_in_0_bits_inputValue_3_tag,
  output        io_out_valid,
  output [3:0]  io_out_bits_bank,
  output [5:0]  io_out_bits_address,
  output [22:0] io_out_bits_inputValue_0_tag,
  output [22:0] io_out_bits_inputValue_1_tag,
  output [22:0] io_out_bits_inputValue_2_tag,
  output [22:0] io_out_bits_inputValue_3_tag
);
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_bank = io_in_0_bits_bank; // @[Arbiter.scala 124:15]
  assign io_out_bits_address = io_in_0_bits_address; // @[Arbiter.scala 124:15]
  assign io_out_bits_inputValue_0_tag = io_in_0_bits_inputValue_0_tag; // @[Arbiter.scala 124:15]
  assign io_out_bits_inputValue_1_tag = io_in_0_bits_inputValue_1_tag; // @[Arbiter.scala 124:15]
  assign io_out_bits_inputValue_2_tag = io_in_0_bits_inputValue_2_tag; // @[Arbiter.scala 124:15]
  assign io_out_bits_inputValue_3_tag = io_in_0_bits_inputValue_3_tag; // @[Arbiter.scala 124:15]
endmodule
module Gem5Cache(
  input         clock,
  input         reset,
  input         io_cpu_0_req_valid,
  input  [31:0] io_cpu_0_req_bits_addr,
  input  [63:0] io_cpu_0_req_bits_data,
  input  [27:0] io_cpu_0_req_bits_command,
  input  [2:0]  io_cpu_0_req_bits_way,
  input  [2:0]  io_cpu_0_req_bits_replaceWay,
  output        io_cpu_0_resp_valid,
  output        io_cpu_0_resp_bits_iswrite,
  output [2:0]  io_cpu_0_resp_bits_way,
  input         io_probe_req_valid,
  input  [31:0] io_probe_req_bits_addr,
  input  [27:0] io_probe_req_bits_command,
  output        io_probe_resp_valid,
  output [2:0]  io_probe_resp_bits_way,
  output        io_probe_multiWay_valid,
  output [2:0]  io_probe_multiWay_bits_way_0,
  output [2:0]  io_probe_multiWay_bits_way_1,
  output [2:0]  io_probe_multiWay_bits_way_2,
  output [2:0]  io_probe_multiWay_bits_way_3,
  output [31:0] io_probe_multiWay_bits_addr,
  input         io_bipassLD_in_valid,
  input  [31:0] io_bipassLD_in_bits_addr,
  input  [3:0]  io_bipassLD_in_bits_way,
  output        io_bipassLD_out_valid,
  output [63:0] io_bipassLD_out_bits_data
);
  wire  biPassModule_clock; // @[AXICache.scala 61:28]
  wire  biPassModule_reset; // @[AXICache.scala 61:28]
  wire  biPassModule_io_in_valid; // @[AXICache.scala 61:28]
  wire [31:0] biPassModule_io_in_bits_addr; // @[AXICache.scala 61:28]
  wire [3:0] biPassModule_io_in_bits_way; // @[AXICache.scala 61:28]
  wire  biPassModule_io_dataMem_in_valid; // @[AXICache.scala 61:28]
  wire [31:0] biPassModule_io_dataMem_in_bits_address; // @[AXICache.scala 61:28]
  wire [63:0] biPassModule_io_dataMem_outputValue_0; // @[AXICache.scala 61:28]
  wire  biPassModule_io_out_valid; // @[AXICache.scala 61:28]
  wire [63:0] biPassModule_io_out_bits_data; // @[AXICache.scala 61:28]
  wire  dataMemory_clock; // @[AXICache.scala 77:26]
  wire  dataMemory_io_read_in_valid; // @[AXICache.scala 77:26]
  wire [31:0] dataMemory_io_read_in_bits_address; // @[AXICache.scala 77:26]
  wire [63:0] dataMemory_io_read_outputValue_0; // @[AXICache.scala 77:26]
  wire  dataMemory_io_write_valid; // @[AXICache.scala 77:26]
  wire [31:0] dataMemory_io_write_bits_address; // @[AXICache.scala 77:26]
  wire [63:0] dataMemory_io_write_bits_inputValue_0; // @[AXICache.scala 77:26]
  wire  metaMemory_clock; // @[AXICache.scala 78:26]
  wire  metaMemory_io_read_in_valid; // @[AXICache.scala 78:26]
  wire [5:0] metaMemory_io_read_in_bits_address; // @[AXICache.scala 78:26]
  wire [22:0] metaMemory_io_read_outputValue_0_tag; // @[AXICache.scala 78:26]
  wire [22:0] metaMemory_io_read_outputValue_1_tag; // @[AXICache.scala 78:26]
  wire [22:0] metaMemory_io_read_outputValue_2_tag; // @[AXICache.scala 78:26]
  wire [22:0] metaMemory_io_read_outputValue_3_tag; // @[AXICache.scala 78:26]
  wire  metaMemory_io_write_valid; // @[AXICache.scala 78:26]
  wire [3:0] metaMemory_io_write_bits_bank; // @[AXICache.scala 78:26]
  wire [5:0] metaMemory_io_write_bits_address; // @[AXICache.scala 78:26]
  wire [22:0] metaMemory_io_write_bits_inputValue_0_tag; // @[AXICache.scala 78:26]
  wire [22:0] metaMemory_io_write_bits_inputValue_1_tag; // @[AXICache.scala 78:26]
  wire [22:0] metaMemory_io_write_bits_inputValue_2_tag; // @[AXICache.scala 78:26]
  wire [22:0] metaMemory_io_write_bits_inputValue_3_tag; // @[AXICache.scala 78:26]
  wire  cacheLogic_0_clock; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_reset; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_cpu_req_ready; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_cpu_req_valid; // @[AXICache.scala 81:28]
  wire [31:0] cacheLogic_0_io_cpu_req_bits_addr; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_0_io_cpu_req_bits_data; // @[AXICache.scala 81:28]
  wire [27:0] cacheLogic_0_io_cpu_req_bits_command; // @[AXICache.scala 81:28]
  wire [2:0] cacheLogic_0_io_cpu_req_bits_way; // @[AXICache.scala 81:28]
  wire [2:0] cacheLogic_0_io_cpu_req_bits_replaceWay; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_cpu_resp_valid; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_cpu_resp_bits_iswrite; // @[AXICache.scala 81:28]
  wire [2:0] cacheLogic_0_io_cpu_resp_bits_way; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_metaMem_write_valid; // @[AXICache.scala 81:28]
  wire [3:0] cacheLogic_0_io_metaMem_write_bits_bank; // @[AXICache.scala 81:28]
  wire [5:0] cacheLogic_0_io_metaMem_write_bits_address; // @[AXICache.scala 81:28]
  wire [22:0] cacheLogic_0_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 81:28]
  wire [22:0] cacheLogic_0_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 81:28]
  wire [22:0] cacheLogic_0_io_metaMem_write_bits_inputValue_2_tag; // @[AXICache.scala 81:28]
  wire [22:0] cacheLogic_0_io_metaMem_write_bits_inputValue_3_tag; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_dataMem_write_valid; // @[AXICache.scala 81:28]
  wire [31:0] cacheLogic_0_io_dataMem_write_bits_address; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_0_io_dataMem_write_bits_inputValue_0; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_validTagBits_write_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_0_io_validTagBits_write_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_validTagBits_write_bits_value; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_validTagBits_read_in_valid; // @[AXICache.scala 81:28]
  wire [63:0] cacheLogic_0_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_validTagBits_read_out_0; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_validTagBits_read_out_1; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_validTagBits_read_out_2; // @[AXICache.scala 81:28]
  wire  cacheLogic_0_io_validTagBits_read_out_3; // @[AXICache.scala 81:28]
  wire  probeUnit_clock; // @[AXICache.scala 85:26]
  wire  probeUnit_reset; // @[AXICache.scala 85:26]
  wire  probeUnit_io_cpu_req_ready; // @[AXICache.scala 85:26]
  wire  probeUnit_io_cpu_req_valid; // @[AXICache.scala 85:26]
  wire [31:0] probeUnit_io_cpu_req_bits_addr; // @[AXICache.scala 85:26]
  wire [27:0] probeUnit_io_cpu_req_bits_command; // @[AXICache.scala 85:26]
  wire  probeUnit_io_cpu_resp_valid; // @[AXICache.scala 85:26]
  wire [2:0] probeUnit_io_cpu_resp_bits_way; // @[AXICache.scala 85:26]
  wire  probeUnit_io_cpu_multiWay_valid; // @[AXICache.scala 85:26]
  wire [2:0] probeUnit_io_cpu_multiWay_bits_way_0; // @[AXICache.scala 85:26]
  wire [2:0] probeUnit_io_cpu_multiWay_bits_way_1; // @[AXICache.scala 85:26]
  wire [2:0] probeUnit_io_cpu_multiWay_bits_way_2; // @[AXICache.scala 85:26]
  wire [2:0] probeUnit_io_cpu_multiWay_bits_way_3; // @[AXICache.scala 85:26]
  wire [31:0] probeUnit_io_cpu_multiWay_bits_addr; // @[AXICache.scala 85:26]
  wire  probeUnit_io_metaMem_read_in_valid; // @[AXICache.scala 85:26]
  wire [5:0] probeUnit_io_metaMem_read_in_bits_address; // @[AXICache.scala 85:26]
  wire [22:0] probeUnit_io_metaMem_read_outputValue_0_tag; // @[AXICache.scala 85:26]
  wire [22:0] probeUnit_io_metaMem_read_outputValue_1_tag; // @[AXICache.scala 85:26]
  wire [22:0] probeUnit_io_metaMem_read_outputValue_2_tag; // @[AXICache.scala 85:26]
  wire [22:0] probeUnit_io_metaMem_read_outputValue_3_tag; // @[AXICache.scala 85:26]
  wire  probeUnit_io_validTagBits_write_valid; // @[AXICache.scala 85:26]
  wire [63:0] probeUnit_io_validTagBits_write_bits_addr; // @[AXICache.scala 85:26]
  wire  probeUnit_io_validTagBits_write_bits_value; // @[AXICache.scala 85:26]
  wire  probeUnit_io_validTagBits_read_in_valid; // @[AXICache.scala 85:26]
  wire [63:0] probeUnit_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 85:26]
  wire  probeUnit_io_validTagBits_read_out_0; // @[AXICache.scala 85:26]
  wire  probeUnit_io_validTagBits_read_out_1; // @[AXICache.scala 85:26]
  wire  probeUnit_io_validTagBits_read_out_2; // @[AXICache.scala 85:26]
  wire  probeUnit_io_validTagBits_read_out_3; // @[AXICache.scala 85:26]
  wire  validTagBits_clock; // @[AXICache.scala 88:28]
  wire  validTagBits_reset; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_0_write_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_0_write_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_0_write_bits_value; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_0_read_in_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_0_read_in_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_0_read_out_0; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_0_read_out_1; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_0_read_out_2; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_0_read_out_3; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_1_write_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_1_write_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_1_write_bits_value; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_1_read_in_valid; // @[AXICache.scala 88:28]
  wire [63:0] validTagBits_io_port_1_read_in_bits_addr; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_1_read_out_0; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_1_read_out_1; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_1_read_out_2; // @[AXICache.scala 88:28]
  wire  validTagBits_io_port_1_read_out_3; // @[AXICache.scala 88:28]
  wire  metaWrArb_io_in_0_valid; // @[AXICache.scala 91:27]
  wire [3:0] metaWrArb_io_in_0_bits_bank; // @[AXICache.scala 91:27]
  wire [5:0] metaWrArb_io_in_0_bits_address; // @[AXICache.scala 91:27]
  wire [22:0] metaWrArb_io_in_0_bits_inputValue_0_tag; // @[AXICache.scala 91:27]
  wire [22:0] metaWrArb_io_in_0_bits_inputValue_1_tag; // @[AXICache.scala 91:27]
  wire [22:0] metaWrArb_io_in_0_bits_inputValue_2_tag; // @[AXICache.scala 91:27]
  wire [22:0] metaWrArb_io_in_0_bits_inputValue_3_tag; // @[AXICache.scala 91:27]
  wire  metaWrArb_io_out_valid; // @[AXICache.scala 91:27]
  wire [3:0] metaWrArb_io_out_bits_bank; // @[AXICache.scala 91:27]
  wire [5:0] metaWrArb_io_out_bits_address; // @[AXICache.scala 91:27]
  wire [22:0] metaWrArb_io_out_bits_inputValue_0_tag; // @[AXICache.scala 91:27]
  wire [22:0] metaWrArb_io_out_bits_inputValue_1_tag; // @[AXICache.scala 91:27]
  wire [22:0] metaWrArb_io_out_bits_inputValue_2_tag; // @[AXICache.scala 91:27]
  wire [22:0] metaWrArb_io_out_bits_inputValue_3_tag; // @[AXICache.scala 91:27]
  bipassLD biPassModule ( // @[AXICache.scala 61:28]
    .clock(biPassModule_clock),
    .reset(biPassModule_reset),
    .io_in_valid(biPassModule_io_in_valid),
    .io_in_bits_addr(biPassModule_io_in_bits_addr),
    .io_in_bits_way(biPassModule_io_in_bits_way),
    .io_dataMem_in_valid(biPassModule_io_dataMem_in_valid),
    .io_dataMem_in_bits_address(biPassModule_io_dataMem_in_bits_address),
    .io_dataMem_outputValue_0(biPassModule_io_dataMem_outputValue_0),
    .io_out_valid(biPassModule_io_out_valid),
    .io_out_bits_data(biPassModule_io_out_bits_data)
  );
  MemBank dataMemory ( // @[AXICache.scala 77:26]
    .clock(dataMemory_clock),
    .io_read_in_valid(dataMemory_io_read_in_valid),
    .io_read_in_bits_address(dataMemory_io_read_in_bits_address),
    .io_read_outputValue_0(dataMemory_io_read_outputValue_0),
    .io_write_valid(dataMemory_io_write_valid),
    .io_write_bits_address(dataMemory_io_write_bits_address),
    .io_write_bits_inputValue_0(dataMemory_io_write_bits_inputValue_0)
  );
  MemBank_1 metaMemory ( // @[AXICache.scala 78:26]
    .clock(metaMemory_clock),
    .io_read_in_valid(metaMemory_io_read_in_valid),
    .io_read_in_bits_address(metaMemory_io_read_in_bits_address),
    .io_read_outputValue_0_tag(metaMemory_io_read_outputValue_0_tag),
    .io_read_outputValue_1_tag(metaMemory_io_read_outputValue_1_tag),
    .io_read_outputValue_2_tag(metaMemory_io_read_outputValue_2_tag),
    .io_read_outputValue_3_tag(metaMemory_io_read_outputValue_3_tag),
    .io_write_valid(metaMemory_io_write_valid),
    .io_write_bits_bank(metaMemory_io_write_bits_bank),
    .io_write_bits_address(metaMemory_io_write_bits_address),
    .io_write_bits_inputValue_0_tag(metaMemory_io_write_bits_inputValue_0_tag),
    .io_write_bits_inputValue_1_tag(metaMemory_io_write_bits_inputValue_1_tag),
    .io_write_bits_inputValue_2_tag(metaMemory_io_write_bits_inputValue_2_tag),
    .io_write_bits_inputValue_3_tag(metaMemory_io_write_bits_inputValue_3_tag)
  );
  Gem5CacheLogic cacheLogic_0 ( // @[AXICache.scala 81:28]
    .clock(cacheLogic_0_clock),
    .reset(cacheLogic_0_reset),
    .io_cpu_req_ready(cacheLogic_0_io_cpu_req_ready),
    .io_cpu_req_valid(cacheLogic_0_io_cpu_req_valid),
    .io_cpu_req_bits_addr(cacheLogic_0_io_cpu_req_bits_addr),
    .io_cpu_req_bits_data(cacheLogic_0_io_cpu_req_bits_data),
    .io_cpu_req_bits_command(cacheLogic_0_io_cpu_req_bits_command),
    .io_cpu_req_bits_way(cacheLogic_0_io_cpu_req_bits_way),
    .io_cpu_req_bits_replaceWay(cacheLogic_0_io_cpu_req_bits_replaceWay),
    .io_cpu_resp_valid(cacheLogic_0_io_cpu_resp_valid),
    .io_cpu_resp_bits_iswrite(cacheLogic_0_io_cpu_resp_bits_iswrite),
    .io_cpu_resp_bits_way(cacheLogic_0_io_cpu_resp_bits_way),
    .io_metaMem_write_valid(cacheLogic_0_io_metaMem_write_valid),
    .io_metaMem_write_bits_bank(cacheLogic_0_io_metaMem_write_bits_bank),
    .io_metaMem_write_bits_address(cacheLogic_0_io_metaMem_write_bits_address),
    .io_metaMem_write_bits_inputValue_0_tag(cacheLogic_0_io_metaMem_write_bits_inputValue_0_tag),
    .io_metaMem_write_bits_inputValue_1_tag(cacheLogic_0_io_metaMem_write_bits_inputValue_1_tag),
    .io_metaMem_write_bits_inputValue_2_tag(cacheLogic_0_io_metaMem_write_bits_inputValue_2_tag),
    .io_metaMem_write_bits_inputValue_3_tag(cacheLogic_0_io_metaMem_write_bits_inputValue_3_tag),
    .io_dataMem_write_valid(cacheLogic_0_io_dataMem_write_valid),
    .io_dataMem_write_bits_address(cacheLogic_0_io_dataMem_write_bits_address),
    .io_dataMem_write_bits_inputValue_0(cacheLogic_0_io_dataMem_write_bits_inputValue_0),
    .io_validTagBits_write_valid(cacheLogic_0_io_validTagBits_write_valid),
    .io_validTagBits_write_bits_addr(cacheLogic_0_io_validTagBits_write_bits_addr),
    .io_validTagBits_write_bits_value(cacheLogic_0_io_validTagBits_write_bits_value),
    .io_validTagBits_read_in_valid(cacheLogic_0_io_validTagBits_read_in_valid),
    .io_validTagBits_read_in_bits_addr(cacheLogic_0_io_validTagBits_read_in_bits_addr),
    .io_validTagBits_read_out_0(cacheLogic_0_io_validTagBits_read_out_0),
    .io_validTagBits_read_out_1(cacheLogic_0_io_validTagBits_read_out_1),
    .io_validTagBits_read_out_2(cacheLogic_0_io_validTagBits_read_out_2),
    .io_validTagBits_read_out_3(cacheLogic_0_io_validTagBits_read_out_3)
  );
  ProbeUnit probeUnit ( // @[AXICache.scala 85:26]
    .clock(probeUnit_clock),
    .reset(probeUnit_reset),
    .io_cpu_req_ready(probeUnit_io_cpu_req_ready),
    .io_cpu_req_valid(probeUnit_io_cpu_req_valid),
    .io_cpu_req_bits_addr(probeUnit_io_cpu_req_bits_addr),
    .io_cpu_req_bits_command(probeUnit_io_cpu_req_bits_command),
    .io_cpu_resp_valid(probeUnit_io_cpu_resp_valid),
    .io_cpu_resp_bits_way(probeUnit_io_cpu_resp_bits_way),
    .io_cpu_multiWay_valid(probeUnit_io_cpu_multiWay_valid),
    .io_cpu_multiWay_bits_way_0(probeUnit_io_cpu_multiWay_bits_way_0),
    .io_cpu_multiWay_bits_way_1(probeUnit_io_cpu_multiWay_bits_way_1),
    .io_cpu_multiWay_bits_way_2(probeUnit_io_cpu_multiWay_bits_way_2),
    .io_cpu_multiWay_bits_way_3(probeUnit_io_cpu_multiWay_bits_way_3),
    .io_cpu_multiWay_bits_addr(probeUnit_io_cpu_multiWay_bits_addr),
    .io_metaMem_read_in_valid(probeUnit_io_metaMem_read_in_valid),
    .io_metaMem_read_in_bits_address(probeUnit_io_metaMem_read_in_bits_address),
    .io_metaMem_read_outputValue_0_tag(probeUnit_io_metaMem_read_outputValue_0_tag),
    .io_metaMem_read_outputValue_1_tag(probeUnit_io_metaMem_read_outputValue_1_tag),
    .io_metaMem_read_outputValue_2_tag(probeUnit_io_metaMem_read_outputValue_2_tag),
    .io_metaMem_read_outputValue_3_tag(probeUnit_io_metaMem_read_outputValue_3_tag),
    .io_validTagBits_write_valid(probeUnit_io_validTagBits_write_valid),
    .io_validTagBits_write_bits_addr(probeUnit_io_validTagBits_write_bits_addr),
    .io_validTagBits_write_bits_value(probeUnit_io_validTagBits_write_bits_value),
    .io_validTagBits_read_in_valid(probeUnit_io_validTagBits_read_in_valid),
    .io_validTagBits_read_in_bits_addr(probeUnit_io_validTagBits_read_in_bits_addr),
    .io_validTagBits_read_out_0(probeUnit_io_validTagBits_read_out_0),
    .io_validTagBits_read_out_1(probeUnit_io_validTagBits_read_out_1),
    .io_validTagBits_read_out_2(probeUnit_io_validTagBits_read_out_2),
    .io_validTagBits_read_out_3(probeUnit_io_validTagBits_read_out_3)
  );
  paralReg_1 validTagBits ( // @[AXICache.scala 88:28]
    .clock(validTagBits_clock),
    .reset(validTagBits_reset),
    .io_port_0_write_valid(validTagBits_io_port_0_write_valid),
    .io_port_0_write_bits_addr(validTagBits_io_port_0_write_bits_addr),
    .io_port_0_write_bits_value(validTagBits_io_port_0_write_bits_value),
    .io_port_0_read_in_valid(validTagBits_io_port_0_read_in_valid),
    .io_port_0_read_in_bits_addr(validTagBits_io_port_0_read_in_bits_addr),
    .io_port_0_read_out_0(validTagBits_io_port_0_read_out_0),
    .io_port_0_read_out_1(validTagBits_io_port_0_read_out_1),
    .io_port_0_read_out_2(validTagBits_io_port_0_read_out_2),
    .io_port_0_read_out_3(validTagBits_io_port_0_read_out_3),
    .io_port_1_write_valid(validTagBits_io_port_1_write_valid),
    .io_port_1_write_bits_addr(validTagBits_io_port_1_write_bits_addr),
    .io_port_1_write_bits_value(validTagBits_io_port_1_write_bits_value),
    .io_port_1_read_in_valid(validTagBits_io_port_1_read_in_valid),
    .io_port_1_read_in_bits_addr(validTagBits_io_port_1_read_in_bits_addr),
    .io_port_1_read_out_0(validTagBits_io_port_1_read_out_0),
    .io_port_1_read_out_1(validTagBits_io_port_1_read_out_1),
    .io_port_1_read_out_2(validTagBits_io_port_1_read_out_2),
    .io_port_1_read_out_3(validTagBits_io_port_1_read_out_3)
  );
  Arbiter_2 metaWrArb ( // @[AXICache.scala 91:27]
    .io_in_0_valid(metaWrArb_io_in_0_valid),
    .io_in_0_bits_bank(metaWrArb_io_in_0_bits_bank),
    .io_in_0_bits_address(metaWrArb_io_in_0_bits_address),
    .io_in_0_bits_inputValue_0_tag(metaWrArb_io_in_0_bits_inputValue_0_tag),
    .io_in_0_bits_inputValue_1_tag(metaWrArb_io_in_0_bits_inputValue_1_tag),
    .io_in_0_bits_inputValue_2_tag(metaWrArb_io_in_0_bits_inputValue_2_tag),
    .io_in_0_bits_inputValue_3_tag(metaWrArb_io_in_0_bits_inputValue_3_tag),
    .io_out_valid(metaWrArb_io_out_valid),
    .io_out_bits_bank(metaWrArb_io_out_bits_bank),
    .io_out_bits_address(metaWrArb_io_out_bits_address),
    .io_out_bits_inputValue_0_tag(metaWrArb_io_out_bits_inputValue_0_tag),
    .io_out_bits_inputValue_1_tag(metaWrArb_io_out_bits_inputValue_1_tag),
    .io_out_bits_inputValue_2_tag(metaWrArb_io_out_bits_inputValue_2_tag),
    .io_out_bits_inputValue_3_tag(metaWrArb_io_out_bits_inputValue_3_tag)
  );
  assign io_cpu_0_resp_valid = cacheLogic_0_io_cpu_resp_valid; // @[AXICache.scala 128:20]
  assign io_cpu_0_resp_bits_iswrite = cacheLogic_0_io_cpu_resp_bits_iswrite; // @[AXICache.scala 128:20]
  assign io_cpu_0_resp_bits_way = cacheLogic_0_io_cpu_resp_bits_way; // @[AXICache.scala 128:20]
  assign io_probe_resp_valid = probeUnit_io_cpu_resp_valid; // @[AXICache.scala 133:17]
  assign io_probe_resp_bits_way = probeUnit_io_cpu_resp_bits_way; // @[AXICache.scala 133:17]
  assign io_probe_multiWay_valid = probeUnit_io_cpu_multiWay_valid; // @[AXICache.scala 133:17]
  assign io_probe_multiWay_bits_way_0 = probeUnit_io_cpu_multiWay_bits_way_0; // @[AXICache.scala 133:17]
  assign io_probe_multiWay_bits_way_1 = probeUnit_io_cpu_multiWay_bits_way_1; // @[AXICache.scala 133:17]
  assign io_probe_multiWay_bits_way_2 = probeUnit_io_cpu_multiWay_bits_way_2; // @[AXICache.scala 133:17]
  assign io_probe_multiWay_bits_way_3 = probeUnit_io_cpu_multiWay_bits_way_3; // @[AXICache.scala 133:17]
  assign io_probe_multiWay_bits_addr = probeUnit_io_cpu_multiWay_bits_addr; // @[AXICache.scala 133:17]
  assign io_bipassLD_out_valid = biPassModule_io_out_valid; // @[AXICache.scala 95:23]
  assign io_bipassLD_out_bits_data = biPassModule_io_out_bits_data; // @[AXICache.scala 95:23]
  assign biPassModule_clock = clock;
  assign biPassModule_reset = reset;
  assign biPassModule_io_in_valid = io_bipassLD_in_valid; // @[AXICache.scala 94:23]
  assign biPassModule_io_in_bits_addr = io_bipassLD_in_bits_addr; // @[AXICache.scala 94:23]
  assign biPassModule_io_in_bits_way = io_bipassLD_in_bits_way; // @[AXICache.scala 94:23]
  assign biPassModule_io_dataMem_outputValue_0 = dataMemory_io_read_outputValue_0; // @[AXICache.scala 97:42]
  assign dataMemory_clock = clock;
  assign dataMemory_io_read_in_valid = biPassModule_io_dataMem_in_valid; // @[AXICache.scala 97:42]
  assign dataMemory_io_read_in_bits_address = biPassModule_io_dataMem_in_bits_address; // @[AXICache.scala 97:42]
  assign dataMemory_io_write_valid = cacheLogic_0_io_dataMem_write_valid; // @[AXICache.scala 104:35]
  assign dataMemory_io_write_bits_address = cacheLogic_0_io_dataMem_write_bits_address; // @[AXICache.scala 104:35]
  assign dataMemory_io_write_bits_inputValue_0 = cacheLogic_0_io_dataMem_write_bits_inputValue_0; // @[AXICache.scala 104:35]
  assign metaMemory_clock = clock;
  assign metaMemory_io_read_in_valid = probeUnit_io_metaMem_read_in_valid; // @[AXICache.scala 98:29]
  assign metaMemory_io_read_in_bits_address = probeUnit_io_metaMem_read_in_bits_address; // @[AXICache.scala 98:29]
  assign metaMemory_io_write_valid = metaWrArb_io_out_valid; // @[AXICache.scala 116:29]
  assign metaMemory_io_write_bits_bank = metaWrArb_io_out_bits_bank; // @[AXICache.scala 113:36]
  assign metaMemory_io_write_bits_address = metaWrArb_io_out_bits_address; // @[AXICache.scala 114:39]
  assign metaMemory_io_write_bits_inputValue_0_tag = metaWrArb_io_out_bits_inputValue_0_tag; // @[AXICache.scala 115:39]
  assign metaMemory_io_write_bits_inputValue_1_tag = metaWrArb_io_out_bits_inputValue_1_tag; // @[AXICache.scala 115:39]
  assign metaMemory_io_write_bits_inputValue_2_tag = metaWrArb_io_out_bits_inputValue_2_tag; // @[AXICache.scala 115:39]
  assign metaMemory_io_write_bits_inputValue_3_tag = metaWrArb_io_out_bits_inputValue_3_tag; // @[AXICache.scala 115:39]
  assign cacheLogic_0_clock = clock;
  assign cacheLogic_0_reset = reset;
  assign cacheLogic_0_io_cpu_req_valid = io_cpu_0_req_valid; // @[AXICache.scala 128:20]
  assign cacheLogic_0_io_cpu_req_bits_addr = io_cpu_0_req_bits_addr; // @[AXICache.scala 128:20]
  assign cacheLogic_0_io_cpu_req_bits_data = io_cpu_0_req_bits_data; // @[AXICache.scala 128:20]
  assign cacheLogic_0_io_cpu_req_bits_command = io_cpu_0_req_bits_command; // @[AXICache.scala 128:20]
  assign cacheLogic_0_io_cpu_req_bits_way = io_cpu_0_req_bits_way; // @[AXICache.scala 128:20]
  assign cacheLogic_0_io_cpu_req_bits_replaceWay = io_cpu_0_req_bits_replaceWay; // @[AXICache.scala 128:20]
  assign cacheLogic_0_io_validTagBits_read_out_0 = validTagBits_io_port_0_read_out_0; // @[AXICache.scala 127:35]
  assign cacheLogic_0_io_validTagBits_read_out_1 = validTagBits_io_port_0_read_out_1; // @[AXICache.scala 127:35]
  assign cacheLogic_0_io_validTagBits_read_out_2 = validTagBits_io_port_0_read_out_2; // @[AXICache.scala 127:35]
  assign cacheLogic_0_io_validTagBits_read_out_3 = validTagBits_io_port_0_read_out_3; // @[AXICache.scala 127:35]
  assign probeUnit_clock = clock;
  assign probeUnit_reset = reset;
  assign probeUnit_io_cpu_req_valid = io_probe_req_valid; // @[AXICache.scala 133:17]
  assign probeUnit_io_cpu_req_bits_addr = io_probe_req_bits_addr; // @[AXICache.scala 133:17]
  assign probeUnit_io_cpu_req_bits_command = io_probe_req_bits_command; // @[AXICache.scala 133:17]
  assign probeUnit_io_metaMem_read_outputValue_0_tag = metaMemory_io_read_outputValue_0_tag; // @[AXICache.scala 98:29]
  assign probeUnit_io_metaMem_read_outputValue_1_tag = metaMemory_io_read_outputValue_1_tag; // @[AXICache.scala 98:29]
  assign probeUnit_io_metaMem_read_outputValue_2_tag = metaMemory_io_read_outputValue_2_tag; // @[AXICache.scala 98:29]
  assign probeUnit_io_metaMem_read_outputValue_3_tag = metaMemory_io_read_outputValue_3_tag; // @[AXICache.scala 98:29]
  assign probeUnit_io_validTagBits_read_out_0 = validTagBits_io_port_1_read_out_0; // @[AXICache.scala 132:29]
  assign probeUnit_io_validTagBits_read_out_1 = validTagBits_io_port_1_read_out_1; // @[AXICache.scala 132:29]
  assign probeUnit_io_validTagBits_read_out_2 = validTagBits_io_port_1_read_out_2; // @[AXICache.scala 132:29]
  assign probeUnit_io_validTagBits_read_out_3 = validTagBits_io_port_1_read_out_3; // @[AXICache.scala 132:29]
  assign validTagBits_clock = clock;
  assign validTagBits_reset = reset;
  assign validTagBits_io_port_0_write_valid = cacheLogic_0_io_validTagBits_write_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_0_write_bits_addr = cacheLogic_0_io_validTagBits_write_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_0_write_bits_value = cacheLogic_0_io_validTagBits_write_bits_value; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_0_read_in_valid = cacheLogic_0_io_validTagBits_read_in_valid; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_0_read_in_bits_addr = cacheLogic_0_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 127:35]
  assign validTagBits_io_port_1_write_valid = probeUnit_io_validTagBits_write_valid; // @[AXICache.scala 132:29]
  assign validTagBits_io_port_1_write_bits_addr = probeUnit_io_validTagBits_write_bits_addr; // @[AXICache.scala 132:29]
  assign validTagBits_io_port_1_write_bits_value = probeUnit_io_validTagBits_write_bits_value; // @[AXICache.scala 132:29]
  assign validTagBits_io_port_1_read_in_valid = probeUnit_io_validTagBits_read_in_valid; // @[AXICache.scala 132:29]
  assign validTagBits_io_port_1_read_in_bits_addr = probeUnit_io_validTagBits_read_in_bits_addr; // @[AXICache.scala 132:29]
  assign metaWrArb_io_in_0_valid = cacheLogic_0_io_metaMem_write_valid; // @[AXICache.scala 108:33]
  assign metaWrArb_io_in_0_bits_bank = cacheLogic_0_io_metaMem_write_bits_bank; // @[AXICache.scala 105:43]
  assign metaWrArb_io_in_0_bits_address = cacheLogic_0_io_metaMem_write_bits_address; // @[AXICache.scala 106:43]
  assign metaWrArb_io_in_0_bits_inputValue_0_tag = cacheLogic_0_io_metaMem_write_bits_inputValue_0_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_0_bits_inputValue_1_tag = cacheLogic_0_io_metaMem_write_bits_inputValue_1_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_0_bits_inputValue_2_tag = cacheLogic_0_io_metaMem_write_bits_inputValue_2_tag; // @[AXICache.scala 107:43]
  assign metaWrArb_io_in_0_bits_inputValue_3_tag = cacheLogic_0_io_metaMem_write_bits_inputValue_3_tag; // @[AXICache.scala 107:43]
endmodule
module FindEmptyLine_2(
  input        io_data_0,
  input        io_data_1,
  input        io_data_2,
  input        io_data_3,
  input        io_data_4,
  input        io_data_5,
  input        io_data_6,
  input        io_data_7,
  output [2:0] io_value_bits
);
  wire  _T = ~io_data_0; // @[elements.scala 74:53]
  wire  _T_1 = ~io_data_1; // @[elements.scala 74:53]
  wire  _T_2 = ~io_data_2; // @[elements.scala 74:53]
  wire  _T_3 = ~io_data_3; // @[elements.scala 74:53]
  wire  _T_4 = ~io_data_4; // @[elements.scala 74:53]
  wire  _T_5 = ~io_data_5; // @[elements.scala 74:53]
  wire  _T_6 = ~io_data_6; // @[elements.scala 74:53]
  wire  _T_7 = ~io_data_7; // @[elements.scala 74:53]
  wire [3:0] _GEN_0 = _T_7 ? 4'h7 : 4'h8; // @[elements.scala 74:66]
  wire [3:0] _GEN_2 = _T_6 ? 4'h6 : _GEN_0; // @[elements.scala 74:66]
  wire [3:0] _GEN_4 = _T_5 ? 4'h5 : _GEN_2; // @[elements.scala 74:66]
  wire [3:0] _GEN_6 = _T_4 ? 4'h4 : _GEN_4; // @[elements.scala 74:66]
  wire [3:0] _GEN_8 = _T_3 ? 4'h3 : _GEN_6; // @[elements.scala 74:66]
  wire [3:0] _GEN_10 = _T_2 ? 4'h2 : _GEN_8; // @[elements.scala 74:66]
  wire [3:0] _GEN_12 = _T_1 ? 4'h1 : _GEN_10; // @[elements.scala 74:66]
  wire [3:0] idx = _T ? 4'h0 : _GEN_12; // @[elements.scala 74:66]
  assign io_value_bits = idx[2:0]; // @[elements.scala 79:19]
endmodule
module Find_2(
  input  [31:0] io_key,
  input  [31:0] io_data_0,
  input  [31:0] io_data_1,
  input  [31:0] io_data_2,
  input  [31:0] io_data_3,
  input  [31:0] io_data_4,
  input  [31:0] io_data_5,
  input  [31:0] io_data_6,
  input  [31:0] io_data_7,
  input         io_valid_0,
  input         io_valid_1,
  input         io_valid_2,
  input         io_valid_3,
  input         io_valid_4,
  input         io_valid_5,
  input         io_valid_6,
  input         io_valid_7,
  output        io_value_valid,
  output [2:0]  io_value_bits
);
  wire  _T = io_data_0 == io_key; // @[elements.scala 35:54]
  wire  _T_1 = io_data_1 == io_key; // @[elements.scala 35:54]
  wire  _T_2 = io_data_2 == io_key; // @[elements.scala 35:54]
  wire  _T_3 = io_data_3 == io_key; // @[elements.scala 35:54]
  wire  _T_4 = io_data_4 == io_key; // @[elements.scala 35:54]
  wire  _T_5 = io_data_5 == io_key; // @[elements.scala 35:54]
  wire  _T_6 = io_data_6 == io_key; // @[elements.scala 35:54]
  wire  _T_7 = io_data_7 == io_key; // @[elements.scala 35:54]
  wire [7:0] bitmap = {_T_7,_T_6,_T_5,_T_4,_T_3,_T_2,_T_1,_T}; // @[Cat.scala 29:58]
  wire [7:0] _T_21 = {io_valid_7,io_valid_6,io_valid_5,io_valid_4,io_valid_3,io_valid_2,io_valid_1,io_valid_0}; // @[elements.scala 36:46]
  wire [7:0] _T_22 = bitmap & _T_21; // @[elements.scala 36:29]
  wire  _T_25 = |_T_22[7:4]; // @[OneHot.scala 32:14]
  wire [3:0] _T_26 = _T_22[7:4] | _T_22[3:0]; // @[OneHot.scala 32:28]
  wire  _T_29 = |_T_26[3:2]; // @[OneHot.scala 32:14]
  wire [1:0] _T_30 = _T_26[3:2] | _T_26[1:0]; // @[OneHot.scala 32:28]
  wire [1:0] _T_32 = {_T_29,_T_30[1]}; // @[Cat.scala 29:58]
  assign io_value_valid = _T_22 != 8'h0; // @[elements.scala 39:20]
  assign io_value_bits = {_T_25,_T_32}; // @[elements.scala 38:19]
endmodule
module TBETable(
  input         clock,
  input         reset,
  input         io_write_0_valid,
  input  [63:0] io_write_0_bits_addr,
  input  [1:0]  io_write_0_bits_command,
  input         io_write_0_bits_mask,
  input  [1:0]  io_write_0_bits_inputTBE_state_state,
  input  [3:0]  io_write_0_bits_inputTBE_way,
  input  [31:0] io_write_0_bits_inputTBE_fields_0,
  input         io_read_valid,
  input  [63:0] io_read_bits_addr,
  output [1:0]  io_outputTBE_bits_state_state,
  output [3:0]  io_outputTBE_bits_way,
  output [31:0] io_outputTBE_bits_fields_0,
  output        io_isFull
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
`endif // RANDOMIZE_REG_INIT
  wire  allocLine_io_data_0; // @[TBE.scala 79:25]
  wire  allocLine_io_data_1; // @[TBE.scala 79:25]
  wire  allocLine_io_data_2; // @[TBE.scala 79:25]
  wire  allocLine_io_data_3; // @[TBE.scala 79:25]
  wire  allocLine_io_data_4; // @[TBE.scala 79:25]
  wire  allocLine_io_data_5; // @[TBE.scala 79:25]
  wire  allocLine_io_data_6; // @[TBE.scala 79:25]
  wire  allocLine_io_data_7; // @[TBE.scala 79:25]
  wire [2:0] allocLine_io_value_bits; // @[TBE.scala 79:25]
  wire [31:0] finder_0_io_key; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_0; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_1; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_2; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_3; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_4; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_5; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_6; // @[TBE.scala 84:24]
  wire [31:0] finder_0_io_data_7; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_0; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_1; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_2; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_3; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_4; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_5; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_6; // @[TBE.scala 84:24]
  wire  finder_0_io_valid_7; // @[TBE.scala 84:24]
  wire  finder_0_io_value_valid; // @[TBE.scala 84:24]
  wire [2:0] finder_0_io_value_bits; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_key; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_0; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_1; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_2; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_3; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_4; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_5; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_6; // @[TBE.scala 84:24]
  wire [31:0] finder_1_io_data_7; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_0; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_1; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_2; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_3; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_4; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_5; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_6; // @[TBE.scala 84:24]
  wire  finder_1_io_valid_7; // @[TBE.scala 84:24]
  wire  finder_1_io_value_valid; // @[TBE.scala 84:24]
  wire [2:0] finder_1_io_value_bits; // @[TBE.scala 84:24]
  reg [1:0] TBEMemory_0_state_state; // @[TBE.scala 62:26]
  reg [3:0] TBEMemory_0_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_0_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_1_state_state; // @[TBE.scala 62:26]
  reg [3:0] TBEMemory_1_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_1_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_2_state_state; // @[TBE.scala 62:26]
  reg [3:0] TBEMemory_2_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_2_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_3_state_state; // @[TBE.scala 62:26]
  reg [3:0] TBEMemory_3_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_3_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_4_state_state; // @[TBE.scala 62:26]
  reg [3:0] TBEMemory_4_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_4_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_5_state_state; // @[TBE.scala 62:26]
  reg [3:0] TBEMemory_5_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_5_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_6_state_state; // @[TBE.scala 62:26]
  reg [3:0] TBEMemory_6_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_6_fields_0; // @[TBE.scala 62:26]
  reg [1:0] TBEMemory_7_state_state; // @[TBE.scala 62:26]
  reg [3:0] TBEMemory_7_way; // @[TBE.scala 62:26]
  reg [31:0] TBEMemory_7_fields_0; // @[TBE.scala 62:26]
  reg  TBEValid_0; // @[TBE.scala 63:25]
  reg  TBEValid_1; // @[TBE.scala 63:25]
  reg  TBEValid_2; // @[TBE.scala 63:25]
  reg  TBEValid_3; // @[TBE.scala 63:25]
  reg  TBEValid_4; // @[TBE.scala 63:25]
  reg  TBEValid_5; // @[TBE.scala 63:25]
  reg  TBEValid_6; // @[TBE.scala 63:25]
  reg  TBEValid_7; // @[TBE.scala 63:25]
  reg [31:0] TBEAddr_0; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_1; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_2; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_3; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_4; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_5; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_6; // @[TBE.scala 64:24]
  reg [31:0] TBEAddr_7; // @[TBE.scala 64:24]
  reg [4:0] counter; // @[TBE.scala 75:24]
  wire [3:0] _T_38 = 4'h8 - 4'h3; // @[TBE.scala 90:40]
  wire [4:0] _GEN_282 = {{1'd0}, _T_38}; // @[TBE.scala 90:26]
  wire  _T_39 = counter > _GEN_282; // @[TBE.scala 90:26]
  wire  _T_40 = _T_39 & io_read_valid; // @[TBE.scala 90:58]
  wire  _T_41 = ~finder_1_io_value_valid; // @[TBE.scala 90:69]
  wire  idxReadValid = finder_1_io_value_valid & io_read_valid; // @[TBE.scala 96:50]
  wire [3:0] idxAlloc = {{1'd0}, allocLine_io_value_bits}; // @[TBE.scala 71:22 TBE.scala 81:12]
  wire  _GEN_283 = 3'h0 == idxAlloc[2:0]; // @[TBE.scala 112:26]
  wire  _GEN_32 = _GEN_283 | TBEValid_0; // @[TBE.scala 112:26]
  wire  _GEN_284 = 3'h1 == idxAlloc[2:0]; // @[TBE.scala 112:26]
  wire  _GEN_33 = _GEN_284 | TBEValid_1; // @[TBE.scala 112:26]
  wire  _GEN_285 = 3'h2 == idxAlloc[2:0]; // @[TBE.scala 112:26]
  wire  _GEN_34 = _GEN_285 | TBEValid_2; // @[TBE.scala 112:26]
  wire  _GEN_286 = 3'h3 == idxAlloc[2:0]; // @[TBE.scala 112:26]
  wire  _GEN_35 = _GEN_286 | TBEValid_3; // @[TBE.scala 112:26]
  wire  _GEN_287 = 3'h4 == idxAlloc[2:0]; // @[TBE.scala 112:26]
  wire  _GEN_36 = _GEN_287 | TBEValid_4; // @[TBE.scala 112:26]
  wire  _GEN_288 = 3'h5 == idxAlloc[2:0]; // @[TBE.scala 112:26]
  wire  _GEN_37 = _GEN_288 | TBEValid_5; // @[TBE.scala 112:26]
  wire  _GEN_289 = 3'h6 == idxAlloc[2:0]; // @[TBE.scala 112:26]
  wire  _GEN_38 = _GEN_289 | TBEValid_6; // @[TBE.scala 112:26]
  wire  _GEN_290 = 3'h7 == idxAlloc[2:0]; // @[TBE.scala 112:26]
  wire  _GEN_39 = _GEN_290 | TBEValid_7; // @[TBE.scala 112:26]
  wire [4:0] _T_51 = counter + 5'h1; // @[TBE.scala 113:26]
  wire  _T_74 = io_write_0_bits_command == 2'h2; // @[TBE.scala 137:46]
  wire  isDealloc_0 = _T_74 & io_write_0_valid; // @[TBE.scala 137:58]
  wire  _T_52 = isDealloc_0 & finder_0_io_value_valid; // @[TBE.scala 114:31]
  wire [3:0] idxUpdate_0 = {{1'd0}, finder_0_io_value_bits}; // @[TBE.scala 73:23 TBE.scala 104:18]
  wire [4:0] _T_59 = counter - 5'h1; // @[TBE.scala 118:26]
  wire  _T_76 = io_write_0_bits_command == 2'h3; // @[TBE.scala 138:44]
  wire  isWrite_0 = _T_76 & io_write_0_valid; // @[TBE.scala 138:55]
  wire  _T_60 = isWrite_0 & finder_0_io_value_valid; // @[TBE.scala 119:29]
  wire  _T_61 = ~io_write_0_bits_mask; // @[TBE.scala 120:35]
  wire  _T_65 = ~reset; // @[TBE.scala 122:15]
  wire [31:0] _GEN_93 = 3'h1 == idxUpdate_0[2:0] ? TBEMemory_1_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 122:15]
  wire [31:0] _GEN_96 = 3'h2 == idxUpdate_0[2:0] ? TBEMemory_2_fields_0 : _GEN_93; // @[TBE.scala 122:15]
  wire [31:0] _GEN_99 = 3'h3 == idxUpdate_0[2:0] ? TBEMemory_3_fields_0 : _GEN_96; // @[TBE.scala 122:15]
  wire [31:0] _GEN_102 = 3'h4 == idxUpdate_0[2:0] ? TBEMemory_4_fields_0 : _GEN_99; // @[TBE.scala 122:15]
  wire [31:0] _GEN_105 = 3'h5 == idxUpdate_0[2:0] ? TBEMemory_5_fields_0 : _GEN_102; // @[TBE.scala 122:15]
  wire [31:0] _GEN_108 = 3'h6 == idxUpdate_0[2:0] ? TBEMemory_6_fields_0 : _GEN_105; // @[TBE.scala 122:15]
  wire [31:0] _GEN_111 = 3'h7 == idxUpdate_0[2:0] ? TBEMemory_7_fields_0 : _GEN_108; // @[TBE.scala 122:15]
  wire  _T_72 = io_write_0_bits_command == 2'h1; // @[TBE.scala 136:44]
  wire  isAlloc_0 = _T_72 & io_write_0_valid; // @[TBE.scala 136:54]
  wire [3:0] idxRead = {{1'd0}, finder_1_io_value_bits}; // @[TBE.scala 72:21 TBE.scala 95:11]
  wire [1:0] _GEN_261 = 3'h1 == idxRead[2:0] ? TBEMemory_1_state_state : TBEMemory_0_state_state; // @[TBE.scala 132:27]
  wire [3:0] _GEN_262 = 3'h1 == idxRead[2:0] ? TBEMemory_1_way : TBEMemory_0_way; // @[TBE.scala 132:27]
  wire [31:0] _GEN_263 = 3'h1 == idxRead[2:0] ? TBEMemory_1_fields_0 : TBEMemory_0_fields_0; // @[TBE.scala 132:27]
  wire [1:0] _GEN_264 = 3'h2 == idxRead[2:0] ? TBEMemory_2_state_state : _GEN_261; // @[TBE.scala 132:27]
  wire [3:0] _GEN_265 = 3'h2 == idxRead[2:0] ? TBEMemory_2_way : _GEN_262; // @[TBE.scala 132:27]
  wire [31:0] _GEN_266 = 3'h2 == idxRead[2:0] ? TBEMemory_2_fields_0 : _GEN_263; // @[TBE.scala 132:27]
  wire [1:0] _GEN_267 = 3'h3 == idxRead[2:0] ? TBEMemory_3_state_state : _GEN_264; // @[TBE.scala 132:27]
  wire [3:0] _GEN_268 = 3'h3 == idxRead[2:0] ? TBEMemory_3_way : _GEN_265; // @[TBE.scala 132:27]
  wire [31:0] _GEN_269 = 3'h3 == idxRead[2:0] ? TBEMemory_3_fields_0 : _GEN_266; // @[TBE.scala 132:27]
  wire [1:0] _GEN_270 = 3'h4 == idxRead[2:0] ? TBEMemory_4_state_state : _GEN_267; // @[TBE.scala 132:27]
  wire [3:0] _GEN_271 = 3'h4 == idxRead[2:0] ? TBEMemory_4_way : _GEN_268; // @[TBE.scala 132:27]
  wire [31:0] _GEN_272 = 3'h4 == idxRead[2:0] ? TBEMemory_4_fields_0 : _GEN_269; // @[TBE.scala 132:27]
  wire [1:0] _GEN_273 = 3'h5 == idxRead[2:0] ? TBEMemory_5_state_state : _GEN_270; // @[TBE.scala 132:27]
  wire [3:0] _GEN_274 = 3'h5 == idxRead[2:0] ? TBEMemory_5_way : _GEN_271; // @[TBE.scala 132:27]
  wire [31:0] _GEN_275 = 3'h5 == idxRead[2:0] ? TBEMemory_5_fields_0 : _GEN_272; // @[TBE.scala 132:27]
  wire [1:0] _GEN_276 = 3'h6 == idxRead[2:0] ? TBEMemory_6_state_state : _GEN_273; // @[TBE.scala 132:27]
  wire [3:0] _GEN_277 = 3'h6 == idxRead[2:0] ? TBEMemory_6_way : _GEN_274; // @[TBE.scala 132:27]
  wire [31:0] _GEN_278 = 3'h6 == idxRead[2:0] ? TBEMemory_6_fields_0 : _GEN_275; // @[TBE.scala 132:27]
  wire [1:0] _GEN_279 = 3'h7 == idxRead[2:0] ? TBEMemory_7_state_state : _GEN_276; // @[TBE.scala 132:27]
  wire [3:0] _GEN_280 = 3'h7 == idxRead[2:0] ? TBEMemory_7_way : _GEN_277; // @[TBE.scala 132:27]
  wire [31:0] _GEN_281 = 3'h7 == idxRead[2:0] ? TBEMemory_7_fields_0 : _GEN_278; // @[TBE.scala 132:27]
  wire  _GEN_291 = ~isAlloc_0; // @[TBE.scala 122:15]
  wire  _GEN_292 = ~_T_52; // @[TBE.scala 122:15]
  wire  _GEN_293 = _GEN_291 & _GEN_292; // @[TBE.scala 122:15]
  wire  _GEN_294 = _GEN_293 & _T_60; // @[TBE.scala 122:15]
  wire  _GEN_295 = _GEN_294 & _T_61; // @[TBE.scala 122:15]
  FindEmptyLine_2 allocLine ( // @[TBE.scala 79:25]
    .io_data_0(allocLine_io_data_0),
    .io_data_1(allocLine_io_data_1),
    .io_data_2(allocLine_io_data_2),
    .io_data_3(allocLine_io_data_3),
    .io_data_4(allocLine_io_data_4),
    .io_data_5(allocLine_io_data_5),
    .io_data_6(allocLine_io_data_6),
    .io_data_7(allocLine_io_data_7),
    .io_value_bits(allocLine_io_value_bits)
  );
  Find_2 finder_0 ( // @[TBE.scala 84:24]
    .io_key(finder_0_io_key),
    .io_data_0(finder_0_io_data_0),
    .io_data_1(finder_0_io_data_1),
    .io_data_2(finder_0_io_data_2),
    .io_data_3(finder_0_io_data_3),
    .io_data_4(finder_0_io_data_4),
    .io_data_5(finder_0_io_data_5),
    .io_data_6(finder_0_io_data_6),
    .io_data_7(finder_0_io_data_7),
    .io_valid_0(finder_0_io_valid_0),
    .io_valid_1(finder_0_io_valid_1),
    .io_valid_2(finder_0_io_valid_2),
    .io_valid_3(finder_0_io_valid_3),
    .io_valid_4(finder_0_io_valid_4),
    .io_valid_5(finder_0_io_valid_5),
    .io_valid_6(finder_0_io_valid_6),
    .io_valid_7(finder_0_io_valid_7),
    .io_value_valid(finder_0_io_value_valid),
    .io_value_bits(finder_0_io_value_bits)
  );
  Find_2 finder_1 ( // @[TBE.scala 84:24]
    .io_key(finder_1_io_key),
    .io_data_0(finder_1_io_data_0),
    .io_data_1(finder_1_io_data_1),
    .io_data_2(finder_1_io_data_2),
    .io_data_3(finder_1_io_data_3),
    .io_data_4(finder_1_io_data_4),
    .io_data_5(finder_1_io_data_5),
    .io_data_6(finder_1_io_data_6),
    .io_data_7(finder_1_io_data_7),
    .io_valid_0(finder_1_io_valid_0),
    .io_valid_1(finder_1_io_valid_1),
    .io_valid_2(finder_1_io_valid_2),
    .io_valid_3(finder_1_io_valid_3),
    .io_valid_4(finder_1_io_valid_4),
    .io_valid_5(finder_1_io_valid_5),
    .io_valid_6(finder_1_io_valid_6),
    .io_valid_7(finder_1_io_valid_7),
    .io_value_valid(finder_1_io_value_valid),
    .io_value_bits(finder_1_io_value_bits)
  );
  assign io_outputTBE_bits_state_state = idxReadValid ? _GEN_279 : 2'h0; // @[TBE.scala 132:21]
  assign io_outputTBE_bits_way = idxReadValid ? _GEN_280 : 4'h4; // @[TBE.scala 132:21]
  assign io_outputTBE_bits_fields_0 = idxReadValid ? _GEN_281 : 32'h0; // @[TBE.scala 132:21]
  assign io_isFull = _T_40 & _T_41; // @[TBE.scala 90:13]
  assign allocLine_io_data_0 = TBEValid_0; // @[TBE.scala 80:21]
  assign allocLine_io_data_1 = TBEValid_1; // @[TBE.scala 80:21]
  assign allocLine_io_data_2 = TBEValid_2; // @[TBE.scala 80:21]
  assign allocLine_io_data_3 = TBEValid_3; // @[TBE.scala 80:21]
  assign allocLine_io_data_4 = TBEValid_4; // @[TBE.scala 80:21]
  assign allocLine_io_data_5 = TBEValid_5; // @[TBE.scala 80:21]
  assign allocLine_io_data_6 = TBEValid_6; // @[TBE.scala 80:21]
  assign allocLine_io_data_7 = TBEValid_7; // @[TBE.scala 80:21]
  assign finder_0_io_key = io_write_0_bits_addr[34:3]; // @[TBE.scala 100:22]
  assign finder_0_io_data_0 = TBEAddr_0; // @[TBE.scala 101:23]
  assign finder_0_io_data_1 = TBEAddr_1; // @[TBE.scala 101:23]
  assign finder_0_io_data_2 = TBEAddr_2; // @[TBE.scala 101:23]
  assign finder_0_io_data_3 = TBEAddr_3; // @[TBE.scala 101:23]
  assign finder_0_io_data_4 = TBEAddr_4; // @[TBE.scala 101:23]
  assign finder_0_io_data_5 = TBEAddr_5; // @[TBE.scala 101:23]
  assign finder_0_io_data_6 = TBEAddr_6; // @[TBE.scala 101:23]
  assign finder_0_io_data_7 = TBEAddr_7; // @[TBE.scala 101:23]
  assign finder_0_io_valid_0 = TBEValid_0; // @[TBE.scala 102:24]
  assign finder_0_io_valid_1 = TBEValid_1; // @[TBE.scala 102:24]
  assign finder_0_io_valid_2 = TBEValid_2; // @[TBE.scala 102:24]
  assign finder_0_io_valid_3 = TBEValid_3; // @[TBE.scala 102:24]
  assign finder_0_io_valid_4 = TBEValid_4; // @[TBE.scala 102:24]
  assign finder_0_io_valid_5 = TBEValid_5; // @[TBE.scala 102:24]
  assign finder_0_io_valid_6 = TBEValid_6; // @[TBE.scala 102:24]
  assign finder_0_io_valid_7 = TBEValid_7; // @[TBE.scala 102:24]
  assign finder_1_io_key = io_read_bits_addr[34:3]; // @[TBE.scala 92:25]
  assign finder_1_io_data_0 = TBEAddr_0; // @[TBE.scala 93:26]
  assign finder_1_io_data_1 = TBEAddr_1; // @[TBE.scala 93:26]
  assign finder_1_io_data_2 = TBEAddr_2; // @[TBE.scala 93:26]
  assign finder_1_io_data_3 = TBEAddr_3; // @[TBE.scala 93:26]
  assign finder_1_io_data_4 = TBEAddr_4; // @[TBE.scala 93:26]
  assign finder_1_io_data_5 = TBEAddr_5; // @[TBE.scala 93:26]
  assign finder_1_io_data_6 = TBEAddr_6; // @[TBE.scala 93:26]
  assign finder_1_io_data_7 = TBEAddr_7; // @[TBE.scala 93:26]
  assign finder_1_io_valid_0 = TBEValid_0; // @[TBE.scala 94:27]
  assign finder_1_io_valid_1 = TBEValid_1; // @[TBE.scala 94:27]
  assign finder_1_io_valid_2 = TBEValid_2; // @[TBE.scala 94:27]
  assign finder_1_io_valid_3 = TBEValid_3; // @[TBE.scala 94:27]
  assign finder_1_io_valid_4 = TBEValid_4; // @[TBE.scala 94:27]
  assign finder_1_io_valid_5 = TBEValid_5; // @[TBE.scala 94:27]
  assign finder_1_io_valid_6 = TBEValid_6; // @[TBE.scala 94:27]
  assign finder_1_io_valid_7 = TBEValid_7; // @[TBE.scala 94:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  TBEMemory_0_state_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  TBEMemory_0_way = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  TBEMemory_0_fields_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  TBEMemory_1_state_state = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  TBEMemory_1_way = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  TBEMemory_1_fields_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  TBEMemory_2_state_state = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  TBEMemory_2_way = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  TBEMemory_2_fields_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  TBEMemory_3_state_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  TBEMemory_3_way = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  TBEMemory_3_fields_0 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  TBEMemory_4_state_state = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  TBEMemory_4_way = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  TBEMemory_4_fields_0 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  TBEMemory_5_state_state = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  TBEMemory_5_way = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  TBEMemory_5_fields_0 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  TBEMemory_6_state_state = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  TBEMemory_6_way = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  TBEMemory_6_fields_0 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  TBEMemory_7_state_state = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  TBEMemory_7_way = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  TBEMemory_7_fields_0 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  TBEValid_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  TBEValid_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  TBEValid_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  TBEValid_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  TBEValid_4 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  TBEValid_5 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  TBEValid_6 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  TBEValid_7 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  TBEAddr_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  TBEAddr_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  TBEAddr_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  TBEAddr_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  TBEAddr_4 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  TBEAddr_5 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  TBEAddr_6 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  TBEAddr_7 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  counter = _RAND_40[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      TBEMemory_0_state_state <= 2'h0;
    end else if (isAlloc_0) begin
      if (3'h0 == idxAlloc[2:0]) begin
        TBEMemory_0_state_state <= io_write_0_bits_inputTBE_state_state;
      end
    end else if (_T_52) begin
      if (3'h0 == idxUpdate_0[2:0]) begin
        TBEMemory_0_state_state <= 2'h0;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h0 == idxUpdate_0[2:0]) begin
          TBEMemory_0_state_state <= io_write_0_bits_inputTBE_state_state;
        end
      end
    end
    if (reset) begin
      TBEMemory_0_way <= 4'h4;
    end else if (isAlloc_0) begin
      if (3'h0 == idxAlloc[2:0]) begin
        TBEMemory_0_way <= io_write_0_bits_inputTBE_way;
      end
    end else if (_T_52) begin
      if (3'h0 == idxUpdate_0[2:0]) begin
        TBEMemory_0_way <= 4'h4;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h0 == idxUpdate_0[2:0]) begin
          TBEMemory_0_way <= io_write_0_bits_inputTBE_way;
        end
      end
    end
    if (reset) begin
      TBEMemory_0_fields_0 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h0 == idxAlloc[2:0]) begin
        TBEMemory_0_fields_0 <= io_write_0_bits_inputTBE_fields_0;
      end
    end else if (_T_52) begin
      if (3'h0 == idxUpdate_0[2:0]) begin
        TBEMemory_0_fields_0 <= 32'h0;
      end
    end else if (_T_60) begin
      if (_T_61) begin
        if (3'h0 == idxUpdate_0[2:0]) begin
          TBEMemory_0_fields_0 <= io_write_0_bits_inputTBE_fields_0;
        end
      end
    end
    if (reset) begin
      TBEMemory_1_state_state <= 2'h0;
    end else if (isAlloc_0) begin
      if (3'h1 == idxAlloc[2:0]) begin
        TBEMemory_1_state_state <= io_write_0_bits_inputTBE_state_state;
      end
    end else if (_T_52) begin
      if (3'h1 == idxUpdate_0[2:0]) begin
        TBEMemory_1_state_state <= 2'h0;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h1 == idxUpdate_0[2:0]) begin
          TBEMemory_1_state_state <= io_write_0_bits_inputTBE_state_state;
        end
      end
    end
    if (reset) begin
      TBEMemory_1_way <= 4'h4;
    end else if (isAlloc_0) begin
      if (3'h1 == idxAlloc[2:0]) begin
        TBEMemory_1_way <= io_write_0_bits_inputTBE_way;
      end
    end else if (_T_52) begin
      if (3'h1 == idxUpdate_0[2:0]) begin
        TBEMemory_1_way <= 4'h4;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h1 == idxUpdate_0[2:0]) begin
          TBEMemory_1_way <= io_write_0_bits_inputTBE_way;
        end
      end
    end
    if (reset) begin
      TBEMemory_1_fields_0 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h1 == idxAlloc[2:0]) begin
        TBEMemory_1_fields_0 <= io_write_0_bits_inputTBE_fields_0;
      end
    end else if (_T_52) begin
      if (3'h1 == idxUpdate_0[2:0]) begin
        TBEMemory_1_fields_0 <= 32'h0;
      end
    end else if (_T_60) begin
      if (_T_61) begin
        if (3'h1 == idxUpdate_0[2:0]) begin
          TBEMemory_1_fields_0 <= io_write_0_bits_inputTBE_fields_0;
        end
      end
    end
    if (reset) begin
      TBEMemory_2_state_state <= 2'h0;
    end else if (isAlloc_0) begin
      if (3'h2 == idxAlloc[2:0]) begin
        TBEMemory_2_state_state <= io_write_0_bits_inputTBE_state_state;
      end
    end else if (_T_52) begin
      if (3'h2 == idxUpdate_0[2:0]) begin
        TBEMemory_2_state_state <= 2'h0;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h2 == idxUpdate_0[2:0]) begin
          TBEMemory_2_state_state <= io_write_0_bits_inputTBE_state_state;
        end
      end
    end
    if (reset) begin
      TBEMemory_2_way <= 4'h4;
    end else if (isAlloc_0) begin
      if (3'h2 == idxAlloc[2:0]) begin
        TBEMemory_2_way <= io_write_0_bits_inputTBE_way;
      end
    end else if (_T_52) begin
      if (3'h2 == idxUpdate_0[2:0]) begin
        TBEMemory_2_way <= 4'h4;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h2 == idxUpdate_0[2:0]) begin
          TBEMemory_2_way <= io_write_0_bits_inputTBE_way;
        end
      end
    end
    if (reset) begin
      TBEMemory_2_fields_0 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h2 == idxAlloc[2:0]) begin
        TBEMemory_2_fields_0 <= io_write_0_bits_inputTBE_fields_0;
      end
    end else if (_T_52) begin
      if (3'h2 == idxUpdate_0[2:0]) begin
        TBEMemory_2_fields_0 <= 32'h0;
      end
    end else if (_T_60) begin
      if (_T_61) begin
        if (3'h2 == idxUpdate_0[2:0]) begin
          TBEMemory_2_fields_0 <= io_write_0_bits_inputTBE_fields_0;
        end
      end
    end
    if (reset) begin
      TBEMemory_3_state_state <= 2'h0;
    end else if (isAlloc_0) begin
      if (3'h3 == idxAlloc[2:0]) begin
        TBEMemory_3_state_state <= io_write_0_bits_inputTBE_state_state;
      end
    end else if (_T_52) begin
      if (3'h3 == idxUpdate_0[2:0]) begin
        TBEMemory_3_state_state <= 2'h0;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h3 == idxUpdate_0[2:0]) begin
          TBEMemory_3_state_state <= io_write_0_bits_inputTBE_state_state;
        end
      end
    end
    if (reset) begin
      TBEMemory_3_way <= 4'h4;
    end else if (isAlloc_0) begin
      if (3'h3 == idxAlloc[2:0]) begin
        TBEMemory_3_way <= io_write_0_bits_inputTBE_way;
      end
    end else if (_T_52) begin
      if (3'h3 == idxUpdate_0[2:0]) begin
        TBEMemory_3_way <= 4'h4;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h3 == idxUpdate_0[2:0]) begin
          TBEMemory_3_way <= io_write_0_bits_inputTBE_way;
        end
      end
    end
    if (reset) begin
      TBEMemory_3_fields_0 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h3 == idxAlloc[2:0]) begin
        TBEMemory_3_fields_0 <= io_write_0_bits_inputTBE_fields_0;
      end
    end else if (_T_52) begin
      if (3'h3 == idxUpdate_0[2:0]) begin
        TBEMemory_3_fields_0 <= 32'h0;
      end
    end else if (_T_60) begin
      if (_T_61) begin
        if (3'h3 == idxUpdate_0[2:0]) begin
          TBEMemory_3_fields_0 <= io_write_0_bits_inputTBE_fields_0;
        end
      end
    end
    if (reset) begin
      TBEMemory_4_state_state <= 2'h0;
    end else if (isAlloc_0) begin
      if (3'h4 == idxAlloc[2:0]) begin
        TBEMemory_4_state_state <= io_write_0_bits_inputTBE_state_state;
      end
    end else if (_T_52) begin
      if (3'h4 == idxUpdate_0[2:0]) begin
        TBEMemory_4_state_state <= 2'h0;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h4 == idxUpdate_0[2:0]) begin
          TBEMemory_4_state_state <= io_write_0_bits_inputTBE_state_state;
        end
      end
    end
    if (reset) begin
      TBEMemory_4_way <= 4'h4;
    end else if (isAlloc_0) begin
      if (3'h4 == idxAlloc[2:0]) begin
        TBEMemory_4_way <= io_write_0_bits_inputTBE_way;
      end
    end else if (_T_52) begin
      if (3'h4 == idxUpdate_0[2:0]) begin
        TBEMemory_4_way <= 4'h4;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h4 == idxUpdate_0[2:0]) begin
          TBEMemory_4_way <= io_write_0_bits_inputTBE_way;
        end
      end
    end
    if (reset) begin
      TBEMemory_4_fields_0 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h4 == idxAlloc[2:0]) begin
        TBEMemory_4_fields_0 <= io_write_0_bits_inputTBE_fields_0;
      end
    end else if (_T_52) begin
      if (3'h4 == idxUpdate_0[2:0]) begin
        TBEMemory_4_fields_0 <= 32'h0;
      end
    end else if (_T_60) begin
      if (_T_61) begin
        if (3'h4 == idxUpdate_0[2:0]) begin
          TBEMemory_4_fields_0 <= io_write_0_bits_inputTBE_fields_0;
        end
      end
    end
    if (reset) begin
      TBEMemory_5_state_state <= 2'h0;
    end else if (isAlloc_0) begin
      if (3'h5 == idxAlloc[2:0]) begin
        TBEMemory_5_state_state <= io_write_0_bits_inputTBE_state_state;
      end
    end else if (_T_52) begin
      if (3'h5 == idxUpdate_0[2:0]) begin
        TBEMemory_5_state_state <= 2'h0;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h5 == idxUpdate_0[2:0]) begin
          TBEMemory_5_state_state <= io_write_0_bits_inputTBE_state_state;
        end
      end
    end
    if (reset) begin
      TBEMemory_5_way <= 4'h4;
    end else if (isAlloc_0) begin
      if (3'h5 == idxAlloc[2:0]) begin
        TBEMemory_5_way <= io_write_0_bits_inputTBE_way;
      end
    end else if (_T_52) begin
      if (3'h5 == idxUpdate_0[2:0]) begin
        TBEMemory_5_way <= 4'h4;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h5 == idxUpdate_0[2:0]) begin
          TBEMemory_5_way <= io_write_0_bits_inputTBE_way;
        end
      end
    end
    if (reset) begin
      TBEMemory_5_fields_0 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h5 == idxAlloc[2:0]) begin
        TBEMemory_5_fields_0 <= io_write_0_bits_inputTBE_fields_0;
      end
    end else if (_T_52) begin
      if (3'h5 == idxUpdate_0[2:0]) begin
        TBEMemory_5_fields_0 <= 32'h0;
      end
    end else if (_T_60) begin
      if (_T_61) begin
        if (3'h5 == idxUpdate_0[2:0]) begin
          TBEMemory_5_fields_0 <= io_write_0_bits_inputTBE_fields_0;
        end
      end
    end
    if (reset) begin
      TBEMemory_6_state_state <= 2'h0;
    end else if (isAlloc_0) begin
      if (3'h6 == idxAlloc[2:0]) begin
        TBEMemory_6_state_state <= io_write_0_bits_inputTBE_state_state;
      end
    end else if (_T_52) begin
      if (3'h6 == idxUpdate_0[2:0]) begin
        TBEMemory_6_state_state <= 2'h0;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h6 == idxUpdate_0[2:0]) begin
          TBEMemory_6_state_state <= io_write_0_bits_inputTBE_state_state;
        end
      end
    end
    if (reset) begin
      TBEMemory_6_way <= 4'h4;
    end else if (isAlloc_0) begin
      if (3'h6 == idxAlloc[2:0]) begin
        TBEMemory_6_way <= io_write_0_bits_inputTBE_way;
      end
    end else if (_T_52) begin
      if (3'h6 == idxUpdate_0[2:0]) begin
        TBEMemory_6_way <= 4'h4;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h6 == idxUpdate_0[2:0]) begin
          TBEMemory_6_way <= io_write_0_bits_inputTBE_way;
        end
      end
    end
    if (reset) begin
      TBEMemory_6_fields_0 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h6 == idxAlloc[2:0]) begin
        TBEMemory_6_fields_0 <= io_write_0_bits_inputTBE_fields_0;
      end
    end else if (_T_52) begin
      if (3'h6 == idxUpdate_0[2:0]) begin
        TBEMemory_6_fields_0 <= 32'h0;
      end
    end else if (_T_60) begin
      if (_T_61) begin
        if (3'h6 == idxUpdate_0[2:0]) begin
          TBEMemory_6_fields_0 <= io_write_0_bits_inputTBE_fields_0;
        end
      end
    end
    if (reset) begin
      TBEMemory_7_state_state <= 2'h0;
    end else if (isAlloc_0) begin
      if (3'h7 == idxAlloc[2:0]) begin
        TBEMemory_7_state_state <= io_write_0_bits_inputTBE_state_state;
      end
    end else if (_T_52) begin
      if (3'h7 == idxUpdate_0[2:0]) begin
        TBEMemory_7_state_state <= 2'h0;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h7 == idxUpdate_0[2:0]) begin
          TBEMemory_7_state_state <= io_write_0_bits_inputTBE_state_state;
        end
      end
    end
    if (reset) begin
      TBEMemory_7_way <= 4'h4;
    end else if (isAlloc_0) begin
      if (3'h7 == idxAlloc[2:0]) begin
        TBEMemory_7_way <= io_write_0_bits_inputTBE_way;
      end
    end else if (_T_52) begin
      if (3'h7 == idxUpdate_0[2:0]) begin
        TBEMemory_7_way <= 4'h4;
      end
    end else if (_T_60) begin
      if (!(_T_61)) begin
        if (3'h7 == idxUpdate_0[2:0]) begin
          TBEMemory_7_way <= io_write_0_bits_inputTBE_way;
        end
      end
    end
    if (reset) begin
      TBEMemory_7_fields_0 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h7 == idxAlloc[2:0]) begin
        TBEMemory_7_fields_0 <= io_write_0_bits_inputTBE_fields_0;
      end
    end else if (_T_52) begin
      if (3'h7 == idxUpdate_0[2:0]) begin
        TBEMemory_7_fields_0 <= 32'h0;
      end
    end else if (_T_60) begin
      if (_T_61) begin
        if (3'h7 == idxUpdate_0[2:0]) begin
          TBEMemory_7_fields_0 <= io_write_0_bits_inputTBE_fields_0;
        end
      end
    end
    if (reset) begin
      TBEValid_0 <= 1'h0;
    end else if (isAlloc_0) begin
      TBEValid_0 <= _GEN_32;
    end else if (_T_52) begin
      if (3'h0 == idxUpdate_0[2:0]) begin
        TBEValid_0 <= 1'h0;
      end
    end
    if (reset) begin
      TBEValid_1 <= 1'h0;
    end else if (isAlloc_0) begin
      TBEValid_1 <= _GEN_33;
    end else if (_T_52) begin
      if (3'h1 == idxUpdate_0[2:0]) begin
        TBEValid_1 <= 1'h0;
      end
    end
    if (reset) begin
      TBEValid_2 <= 1'h0;
    end else if (isAlloc_0) begin
      TBEValid_2 <= _GEN_34;
    end else if (_T_52) begin
      if (3'h2 == idxUpdate_0[2:0]) begin
        TBEValid_2 <= 1'h0;
      end
    end
    if (reset) begin
      TBEValid_3 <= 1'h0;
    end else if (isAlloc_0) begin
      TBEValid_3 <= _GEN_35;
    end else if (_T_52) begin
      if (3'h3 == idxUpdate_0[2:0]) begin
        TBEValid_3 <= 1'h0;
      end
    end
    if (reset) begin
      TBEValid_4 <= 1'h0;
    end else if (isAlloc_0) begin
      TBEValid_4 <= _GEN_36;
    end else if (_T_52) begin
      if (3'h4 == idxUpdate_0[2:0]) begin
        TBEValid_4 <= 1'h0;
      end
    end
    if (reset) begin
      TBEValid_5 <= 1'h0;
    end else if (isAlloc_0) begin
      TBEValid_5 <= _GEN_37;
    end else if (_T_52) begin
      if (3'h5 == idxUpdate_0[2:0]) begin
        TBEValid_5 <= 1'h0;
      end
    end
    if (reset) begin
      TBEValid_6 <= 1'h0;
    end else if (isAlloc_0) begin
      TBEValid_6 <= _GEN_38;
    end else if (_T_52) begin
      if (3'h6 == idxUpdate_0[2:0]) begin
        TBEValid_6 <= 1'h0;
      end
    end
    if (reset) begin
      TBEValid_7 <= 1'h0;
    end else if (isAlloc_0) begin
      TBEValid_7 <= _GEN_39;
    end else if (_T_52) begin
      if (3'h7 == idxUpdate_0[2:0]) begin
        TBEValid_7 <= 1'h0;
      end
    end
    if (reset) begin
      TBEAddr_0 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h0 == idxAlloc[2:0]) begin
        TBEAddr_0 <= io_write_0_bits_addr[34:3];
      end
    end else if (_T_52) begin
      if (3'h0 == idxUpdate_0[2:0]) begin
        TBEAddr_0 <= 32'h0;
      end
    end
    if (reset) begin
      TBEAddr_1 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h1 == idxAlloc[2:0]) begin
        TBEAddr_1 <= io_write_0_bits_addr[34:3];
      end
    end else if (_T_52) begin
      if (3'h1 == idxUpdate_0[2:0]) begin
        TBEAddr_1 <= 32'h0;
      end
    end
    if (reset) begin
      TBEAddr_2 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h2 == idxAlloc[2:0]) begin
        TBEAddr_2 <= io_write_0_bits_addr[34:3];
      end
    end else if (_T_52) begin
      if (3'h2 == idxUpdate_0[2:0]) begin
        TBEAddr_2 <= 32'h0;
      end
    end
    if (reset) begin
      TBEAddr_3 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h3 == idxAlloc[2:0]) begin
        TBEAddr_3 <= io_write_0_bits_addr[34:3];
      end
    end else if (_T_52) begin
      if (3'h3 == idxUpdate_0[2:0]) begin
        TBEAddr_3 <= 32'h0;
      end
    end
    if (reset) begin
      TBEAddr_4 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h4 == idxAlloc[2:0]) begin
        TBEAddr_4 <= io_write_0_bits_addr[34:3];
      end
    end else if (_T_52) begin
      if (3'h4 == idxUpdate_0[2:0]) begin
        TBEAddr_4 <= 32'h0;
      end
    end
    if (reset) begin
      TBEAddr_5 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h5 == idxAlloc[2:0]) begin
        TBEAddr_5 <= io_write_0_bits_addr[34:3];
      end
    end else if (_T_52) begin
      if (3'h5 == idxUpdate_0[2:0]) begin
        TBEAddr_5 <= 32'h0;
      end
    end
    if (reset) begin
      TBEAddr_6 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h6 == idxAlloc[2:0]) begin
        TBEAddr_6 <= io_write_0_bits_addr[34:3];
      end
    end else if (_T_52) begin
      if (3'h6 == idxUpdate_0[2:0]) begin
        TBEAddr_6 <= 32'h0;
      end
    end
    if (reset) begin
      TBEAddr_7 <= 32'h0;
    end else if (isAlloc_0) begin
      if (3'h7 == idxAlloc[2:0]) begin
        TBEAddr_7 <= io_write_0_bits_addr[34:3];
      end
    end else if (_T_52) begin
      if (3'h7 == idxUpdate_0[2:0]) begin
        TBEAddr_7 <= 32'h0;
      end
    end
    if (reset) begin
      counter <= 5'h0;
    end else if (isAlloc_0) begin
      counter <= _T_51;
    end else if (_T_52) begin
      counter <= _T_59;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & _T_65) begin
          $fwrite(32'h80000002,"TBE Field Check %d\n",_GEN_111); // @[TBE.scala 122:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module lockVector(
  input         clock,
  input         reset,
  input         io_lock_in_valid,
  input  [31:0] io_lock_in_bits_addr,
  output        io_probe_out_valid,
  output        io_probe_out_bits,
  input         io_probe_in_valid,
  input  [31:0] io_probe_in_bits_addr,
  input         io_unLock_0_in_valid,
  input  [31:0] io_unLock_0_in_bits_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] finder_0_io_key; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_0; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_1; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_2; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_3; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_4; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_5; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_6; // @[elements.scala 158:28]
  wire [31:0] finder_0_io_data_7; // @[elements.scala 158:28]
  wire  finder_0_io_valid_0; // @[elements.scala 158:28]
  wire  finder_0_io_valid_1; // @[elements.scala 158:28]
  wire  finder_0_io_valid_2; // @[elements.scala 158:28]
  wire  finder_0_io_valid_3; // @[elements.scala 158:28]
  wire  finder_0_io_valid_4; // @[elements.scala 158:28]
  wire  finder_0_io_valid_5; // @[elements.scala 158:28]
  wire  finder_0_io_valid_6; // @[elements.scala 158:28]
  wire  finder_0_io_valid_7; // @[elements.scala 158:28]
  wire  finder_0_io_value_valid; // @[elements.scala 158:28]
  wire [2:0] finder_0_io_value_bits; // @[elements.scala 158:28]
  reg [31:0] addrVec_0; // @[elements.scala 148:26]
  reg [31:0] addrVec_1; // @[elements.scala 148:26]
  reg [31:0] addrVec_2; // @[elements.scala 148:26]
  reg [31:0] addrVec_3; // @[elements.scala 148:26]
  reg [31:0] addrVec_4; // @[elements.scala 148:26]
  reg [31:0] addrVec_5; // @[elements.scala 148:26]
  reg [31:0] addrVec_6; // @[elements.scala 148:26]
  reg [31:0] addrVec_7; // @[elements.scala 148:26]
  reg  valid_0; // @[elements.scala 149:26]
  reg  valid_1; // @[elements.scala 149:26]
  reg  valid_2; // @[elements.scala 149:26]
  reg  valid_3; // @[elements.scala 149:26]
  reg  valid_4; // @[elements.scala 149:26]
  reg  valid_5; // @[elements.scala 149:26]
  reg  valid_6; // @[elements.scala 149:26]
  reg  valid_7; // @[elements.scala 149:26]
  wire [31:0] _GEN_57 = {{3'd0}, io_probe_in_bits_addr[31:3]}; // @[elements.scala 175:53]
  wire  _T_23 = addrVec_7 == _GEN_57; // @[elements.scala 175:53]
  wire  _T_21 = addrVec_6 == _GEN_57; // @[elements.scala 175:53]
  wire  _T_19 = addrVec_5 == _GEN_57; // @[elements.scala 175:53]
  wire  _T_17 = addrVec_4 == _GEN_57; // @[elements.scala 175:53]
  wire  _T_15 = addrVec_3 == _GEN_57; // @[elements.scala 175:53]
  wire  _T_13 = addrVec_2 == _GEN_57; // @[elements.scala 175:53]
  wire  _T_11 = addrVec_1 == _GEN_57; // @[elements.scala 175:53]
  wire  _T_9 = addrVec_0 == _GEN_57; // @[elements.scala 175:53]
  wire [7:0] bitmapProbe = {_T_23,_T_21,_T_19,_T_17,_T_15,_T_13,_T_11,_T_9}; // @[Cat.scala 29:58]
  wire [7:0] _T_69 = {valid_7,valid_6,valid_5,valid_4,valid_3,valid_2,valid_1,valid_0}; // @[elements.scala 201:45]
  wire [7:0] _T_70 = bitmapProbe & _T_69; // @[elements.scala 201:31]
  wire  isLocked = _T_70 != 8'h0; // @[elements.scala 201:49]
  wire  _T_4 = ~isLocked; // @[elements.scala 171:28]
  wire  write = _T_4 & io_lock_in_valid; // @[elements.scala 171:38]
  wire  _T_53 = io_unLock_0_in_valid & finder_0_io_value_valid; // @[elements.scala 189:23]
  wire [7:0] idxUnlock_0 = {{5'd0}, finder_0_io_value_bits}; // @[elements.scala 155:26 elements.scala 185:22]
  wire  _GEN_0 = 3'h0 == idxUnlock_0[2:0] ? 1'h0 : valid_0; // @[elements.scala 190:33]
  wire  _GEN_1 = 3'h1 == idxUnlock_0[2:0] ? 1'h0 : valid_1; // @[elements.scala 190:33]
  wire  _GEN_2 = 3'h2 == idxUnlock_0[2:0] ? 1'h0 : valid_2; // @[elements.scala 190:33]
  wire  _GEN_3 = 3'h3 == idxUnlock_0[2:0] ? 1'h0 : valid_3; // @[elements.scala 190:33]
  wire  _GEN_4 = 3'h4 == idxUnlock_0[2:0] ? 1'h0 : valid_4; // @[elements.scala 190:33]
  wire  _GEN_5 = 3'h5 == idxUnlock_0[2:0] ? 1'h0 : valid_5; // @[elements.scala 190:33]
  wire  _GEN_6 = 3'h6 == idxUnlock_0[2:0] ? 1'h0 : valid_6; // @[elements.scala 190:33]
  wire  _GEN_7 = 3'h7 == idxUnlock_0[2:0] ? 1'h0 : valid_7; // @[elements.scala 190:33]
  wire  _GEN_8 = _T_53 ? _GEN_0 : valid_0; // @[elements.scala 189:52]
  wire  _GEN_9 = _T_53 ? _GEN_1 : valid_1; // @[elements.scala 189:52]
  wire  _GEN_10 = _T_53 ? _GEN_2 : valid_2; // @[elements.scala 189:52]
  wire  _GEN_11 = _T_53 ? _GEN_3 : valid_3; // @[elements.scala 189:52]
  wire  _GEN_12 = _T_53 ? _GEN_4 : valid_4; // @[elements.scala 189:52]
  wire  _GEN_13 = _T_53 ? _GEN_5 : valid_5; // @[elements.scala 189:52]
  wire  _GEN_14 = _T_53 ? _GEN_6 : valid_6; // @[elements.scala 189:52]
  wire  _GEN_15 = _T_53 ? _GEN_7 : valid_7; // @[elements.scala 189:52]
  wire  _T_55 = ~valid_0; // @[elements.scala 196:46]
  wire  _T_56 = ~valid_1; // @[elements.scala 196:46]
  wire  _T_57 = ~valid_2; // @[elements.scala 196:46]
  wire  _T_58 = ~valid_3; // @[elements.scala 196:46]
  wire  _T_59 = ~valid_4; // @[elements.scala 196:46]
  wire  _T_60 = ~valid_5; // @[elements.scala 196:46]
  wire  _T_61 = ~valid_6; // @[elements.scala 196:46]
  wire  _T_62 = ~valid_7; // @[elements.scala 196:46]
  wire [3:0] _GEN_16 = _T_62 ? 4'h7 : 4'h8; // @[elements.scala 196:59]
  wire [3:0] _GEN_17 = _T_61 ? 4'h6 : _GEN_16; // @[elements.scala 196:59]
  wire [3:0] _GEN_18 = _T_60 ? 4'h5 : _GEN_17; // @[elements.scala 196:59]
  wire [3:0] _GEN_19 = _T_59 ? 4'h4 : _GEN_18; // @[elements.scala 196:59]
  wire [3:0] _GEN_20 = _T_58 ? 4'h3 : _GEN_19; // @[elements.scala 196:59]
  wire [3:0] _GEN_21 = _T_57 ? 4'h2 : _GEN_20; // @[elements.scala 196:59]
  wire [3:0] _GEN_22 = _T_56 ? 4'h1 : _GEN_21; // @[elements.scala 196:59]
  wire [3:0] _GEN_23 = _T_55 ? 4'h0 : _GEN_22; // @[elements.scala 196:59]
  wire [7:0] idxLocking = {{4'd0}, _GEN_23}; // @[elements.scala 153:26 elements.scala 177:16 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28 elements.scala 197:28]
  wire [31:0] _addrVec_T_72 = {{3'd0}, io_lock_in_bits_addr[31:3]}; // @[elements.scala 208:29 elements.scala 208:29]
  wire  _GEN_65 = 3'h0 == idxLocking[2:0]; // @[elements.scala 212:27]
  wire  _GEN_41 = _GEN_65 | _GEN_8; // @[elements.scala 212:27]
  wire  _GEN_66 = 3'h1 == idxLocking[2:0]; // @[elements.scala 212:27]
  wire  _GEN_42 = _GEN_66 | _GEN_9; // @[elements.scala 212:27]
  wire  _GEN_67 = 3'h2 == idxLocking[2:0]; // @[elements.scala 212:27]
  wire  _GEN_43 = _GEN_67 | _GEN_10; // @[elements.scala 212:27]
  wire  _GEN_68 = 3'h3 == idxLocking[2:0]; // @[elements.scala 212:27]
  wire  _GEN_44 = _GEN_68 | _GEN_11; // @[elements.scala 212:27]
  wire  _GEN_69 = 3'h4 == idxLocking[2:0]; // @[elements.scala 212:27]
  wire  _GEN_45 = _GEN_69 | _GEN_12; // @[elements.scala 212:27]
  wire  _GEN_70 = 3'h5 == idxLocking[2:0]; // @[elements.scala 212:27]
  wire  _GEN_46 = _GEN_70 | _GEN_13; // @[elements.scala 212:27]
  wire  _GEN_71 = 3'h6 == idxLocking[2:0]; // @[elements.scala 212:27]
  wire  _GEN_47 = _GEN_71 | _GEN_14; // @[elements.scala 212:27]
  wire  _GEN_72 = 3'h7 == idxLocking[2:0]; // @[elements.scala 212:27]
  wire  _GEN_48 = _GEN_72 | _GEN_15; // @[elements.scala 212:27]
  Find_2 finder_0 ( // @[elements.scala 158:28]
    .io_key(finder_0_io_key),
    .io_data_0(finder_0_io_data_0),
    .io_data_1(finder_0_io_data_1),
    .io_data_2(finder_0_io_data_2),
    .io_data_3(finder_0_io_data_3),
    .io_data_4(finder_0_io_data_4),
    .io_data_5(finder_0_io_data_5),
    .io_data_6(finder_0_io_data_6),
    .io_data_7(finder_0_io_data_7),
    .io_valid_0(finder_0_io_valid_0),
    .io_valid_1(finder_0_io_valid_1),
    .io_valid_2(finder_0_io_valid_2),
    .io_valid_3(finder_0_io_valid_3),
    .io_valid_4(finder_0_io_valid_4),
    .io_valid_5(finder_0_io_valid_5),
    .io_valid_6(finder_0_io_valid_6),
    .io_valid_7(finder_0_io_valid_7),
    .io_value_valid(finder_0_io_value_valid),
    .io_value_bits(finder_0_io_value_bits)
  );
  assign io_probe_out_valid = io_probe_in_valid; // @[elements.scala 203:24]
  assign io_probe_out_bits = _T_70 != 8'h0; // @[elements.scala 202:23]
  assign finder_0_io_key = {{3'd0}, io_unLock_0_in_bits_addr[31:3]}; // @[elements.scala 183:26]
  assign finder_0_io_data_0 = addrVec_0; // @[elements.scala 182:27]
  assign finder_0_io_data_1 = addrVec_1; // @[elements.scala 182:27]
  assign finder_0_io_data_2 = addrVec_2; // @[elements.scala 182:27]
  assign finder_0_io_data_3 = addrVec_3; // @[elements.scala 182:27]
  assign finder_0_io_data_4 = addrVec_4; // @[elements.scala 182:27]
  assign finder_0_io_data_5 = addrVec_5; // @[elements.scala 182:27]
  assign finder_0_io_data_6 = addrVec_6; // @[elements.scala 182:27]
  assign finder_0_io_data_7 = addrVec_7; // @[elements.scala 182:27]
  assign finder_0_io_valid_0 = valid_0; // @[elements.scala 184:28]
  assign finder_0_io_valid_1 = valid_1; // @[elements.scala 184:28]
  assign finder_0_io_valid_2 = valid_2; // @[elements.scala 184:28]
  assign finder_0_io_valid_3 = valid_3; // @[elements.scala 184:28]
  assign finder_0_io_valid_4 = valid_4; // @[elements.scala 184:28]
  assign finder_0_io_valid_5 = valid_5; // @[elements.scala 184:28]
  assign finder_0_io_valid_6 = valid_6; // @[elements.scala 184:28]
  assign finder_0_io_valid_7 = valid_7; // @[elements.scala 184:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addrVec_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  addrVec_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  addrVec_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  addrVec_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  addrVec_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  addrVec_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  addrVec_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  addrVec_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  valid_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_4 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_5 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_6 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_7 = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addrVec_0 <= 32'h0;
    end else if (write) begin
      if (3'h0 == idxLocking[2:0]) begin
        addrVec_0 <= _addrVec_T_72;
      end
    end
    if (reset) begin
      addrVec_1 <= 32'h0;
    end else if (write) begin
      if (3'h1 == idxLocking[2:0]) begin
        addrVec_1 <= _addrVec_T_72;
      end
    end
    if (reset) begin
      addrVec_2 <= 32'h0;
    end else if (write) begin
      if (3'h2 == idxLocking[2:0]) begin
        addrVec_2 <= _addrVec_T_72;
      end
    end
    if (reset) begin
      addrVec_3 <= 32'h0;
    end else if (write) begin
      if (3'h3 == idxLocking[2:0]) begin
        addrVec_3 <= _addrVec_T_72;
      end
    end
    if (reset) begin
      addrVec_4 <= 32'h0;
    end else if (write) begin
      if (3'h4 == idxLocking[2:0]) begin
        addrVec_4 <= _addrVec_T_72;
      end
    end
    if (reset) begin
      addrVec_5 <= 32'h0;
    end else if (write) begin
      if (3'h5 == idxLocking[2:0]) begin
        addrVec_5 <= _addrVec_T_72;
      end
    end
    if (reset) begin
      addrVec_6 <= 32'h0;
    end else if (write) begin
      if (3'h6 == idxLocking[2:0]) begin
        addrVec_6 <= _addrVec_T_72;
      end
    end
    if (reset) begin
      addrVec_7 <= 32'h0;
    end else if (write) begin
      if (3'h7 == idxLocking[2:0]) begin
        addrVec_7 <= _addrVec_T_72;
      end
    end
    if (reset) begin
      valid_0 <= 1'h0;
    end else if (write) begin
      valid_0 <= _GEN_41;
    end else if (_T_53) begin
      if (3'h0 == idxUnlock_0[2:0]) begin
        valid_0 <= 1'h0;
      end
    end
    if (reset) begin
      valid_1 <= 1'h0;
    end else if (write) begin
      valid_1 <= _GEN_42;
    end else if (_T_53) begin
      if (3'h1 == idxUnlock_0[2:0]) begin
        valid_1 <= 1'h0;
      end
    end
    if (reset) begin
      valid_2 <= 1'h0;
    end else if (write) begin
      valid_2 <= _GEN_43;
    end else if (_T_53) begin
      if (3'h2 == idxUnlock_0[2:0]) begin
        valid_2 <= 1'h0;
      end
    end
    if (reset) begin
      valid_3 <= 1'h0;
    end else if (write) begin
      valid_3 <= _GEN_44;
    end else if (_T_53) begin
      if (3'h3 == idxUnlock_0[2:0]) begin
        valid_3 <= 1'h0;
      end
    end
    if (reset) begin
      valid_4 <= 1'h0;
    end else if (write) begin
      valid_4 <= _GEN_45;
    end else if (_T_53) begin
      if (3'h4 == idxUnlock_0[2:0]) begin
        valid_4 <= 1'h0;
      end
    end
    if (reset) begin
      valid_5 <= 1'h0;
    end else if (write) begin
      valid_5 <= _GEN_46;
    end else if (_T_53) begin
      if (3'h5 == idxUnlock_0[2:0]) begin
        valid_5 <= 1'h0;
      end
    end
    if (reset) begin
      valid_6 <= 1'h0;
    end else if (write) begin
      valid_6 <= _GEN_47;
    end else if (_T_53) begin
      if (3'h6 == idxUnlock_0[2:0]) begin
        valid_6 <= 1'h0;
      end
    end
    if (reset) begin
      valid_7 <= 1'h0;
    end else if (write) begin
      valid_7 <= _GEN_48;
    end else if (_T_53) begin
      if (3'h7 == idxUnlock_0[2:0]) begin
        valid_7 <= 1'h0;
      end
    end
  end
endmodule
module stateMem(
  input         clock,
  input         reset,
  input         io_in_0_valid,
  input  [1:0]  io_in_0_bits_state_state,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_way,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [2:0]  io_in_1_bits_way,
  output        io_out_valid,
  output [1:0]  io_out_bits_state
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] states_0_state; // @[elements.scala 234:25]
  reg [1:0] states_1_state; // @[elements.scala 234:25]
  reg [1:0] states_2_state; // @[elements.scala 234:25]
  reg [1:0] states_3_state; // @[elements.scala 234:25]
  reg [1:0] states_4_state; // @[elements.scala 234:25]
  reg [1:0] states_5_state; // @[elements.scala 234:25]
  reg [1:0] states_6_state; // @[elements.scala 234:25]
  reg [1:0] states_7_state; // @[elements.scala 234:25]
  reg [1:0] states_8_state; // @[elements.scala 234:25]
  reg [1:0] states_9_state; // @[elements.scala 234:25]
  reg [1:0] states_10_state; // @[elements.scala 234:25]
  reg [1:0] states_11_state; // @[elements.scala 234:25]
  reg [1:0] states_12_state; // @[elements.scala 234:25]
  reg [1:0] states_13_state; // @[elements.scala 234:25]
  reg [1:0] states_14_state; // @[elements.scala 234:25]
  reg [1:0] states_15_state; // @[elements.scala 234:25]
  reg [1:0] states_16_state; // @[elements.scala 234:25]
  reg [1:0] states_17_state; // @[elements.scala 234:25]
  reg [1:0] states_18_state; // @[elements.scala 234:25]
  reg [1:0] states_19_state; // @[elements.scala 234:25]
  reg [1:0] states_20_state; // @[elements.scala 234:25]
  reg [1:0] states_21_state; // @[elements.scala 234:25]
  reg [1:0] states_22_state; // @[elements.scala 234:25]
  reg [1:0] states_23_state; // @[elements.scala 234:25]
  reg [1:0] states_24_state; // @[elements.scala 234:25]
  reg [1:0] states_25_state; // @[elements.scala 234:25]
  reg [1:0] states_26_state; // @[elements.scala 234:25]
  reg [1:0] states_27_state; // @[elements.scala 234:25]
  reg [1:0] states_28_state; // @[elements.scala 234:25]
  reg [1:0] states_29_state; // @[elements.scala 234:25]
  reg [1:0] states_30_state; // @[elements.scala 234:25]
  reg [1:0] states_31_state; // @[elements.scala 234:25]
  reg [1:0] states_32_state; // @[elements.scala 234:25]
  reg [1:0] states_33_state; // @[elements.scala 234:25]
  reg [1:0] states_34_state; // @[elements.scala 234:25]
  reg [1:0] states_35_state; // @[elements.scala 234:25]
  reg [1:0] states_36_state; // @[elements.scala 234:25]
  reg [1:0] states_37_state; // @[elements.scala 234:25]
  reg [1:0] states_38_state; // @[elements.scala 234:25]
  reg [1:0] states_39_state; // @[elements.scala 234:25]
  reg [1:0] states_40_state; // @[elements.scala 234:25]
  reg [1:0] states_41_state; // @[elements.scala 234:25]
  reg [1:0] states_42_state; // @[elements.scala 234:25]
  reg [1:0] states_43_state; // @[elements.scala 234:25]
  reg [1:0] states_44_state; // @[elements.scala 234:25]
  reg [1:0] states_45_state; // @[elements.scala 234:25]
  reg [1:0] states_46_state; // @[elements.scala 234:25]
  reg [1:0] states_47_state; // @[elements.scala 234:25]
  reg [1:0] states_48_state; // @[elements.scala 234:25]
  reg [1:0] states_49_state; // @[elements.scala 234:25]
  reg [1:0] states_50_state; // @[elements.scala 234:25]
  reg [1:0] states_51_state; // @[elements.scala 234:25]
  reg [1:0] states_52_state; // @[elements.scala 234:25]
  reg [1:0] states_53_state; // @[elements.scala 234:25]
  reg [1:0] states_54_state; // @[elements.scala 234:25]
  reg [1:0] states_55_state; // @[elements.scala 234:25]
  reg [1:0] states_56_state; // @[elements.scala 234:25]
  reg [1:0] states_57_state; // @[elements.scala 234:25]
  reg [1:0] states_58_state; // @[elements.scala 234:25]
  reg [1:0] states_59_state; // @[elements.scala 234:25]
  reg [1:0] states_60_state; // @[elements.scala 234:25]
  reg [1:0] states_61_state; // @[elements.scala 234:25]
  reg [1:0] states_62_state; // @[elements.scala 234:25]
  reg [1:0] states_63_state; // @[elements.scala 234:25]
  reg [1:0] states_64_state; // @[elements.scala 234:25]
  reg [1:0] states_65_state; // @[elements.scala 234:25]
  reg [1:0] states_66_state; // @[elements.scala 234:25]
  reg [1:0] states_67_state; // @[elements.scala 234:25]
  reg [1:0] states_68_state; // @[elements.scala 234:25]
  reg [1:0] states_69_state; // @[elements.scala 234:25]
  reg [1:0] states_70_state; // @[elements.scala 234:25]
  reg [1:0] states_71_state; // @[elements.scala 234:25]
  reg [1:0] states_72_state; // @[elements.scala 234:25]
  reg [1:0] states_73_state; // @[elements.scala 234:25]
  reg [1:0] states_74_state; // @[elements.scala 234:25]
  reg [1:0] states_75_state; // @[elements.scala 234:25]
  reg [1:0] states_76_state; // @[elements.scala 234:25]
  reg [1:0] states_77_state; // @[elements.scala 234:25]
  reg [1:0] states_78_state; // @[elements.scala 234:25]
  reg [1:0] states_79_state; // @[elements.scala 234:25]
  reg [1:0] states_80_state; // @[elements.scala 234:25]
  reg [1:0] states_81_state; // @[elements.scala 234:25]
  reg [1:0] states_82_state; // @[elements.scala 234:25]
  reg [1:0] states_83_state; // @[elements.scala 234:25]
  reg [1:0] states_84_state; // @[elements.scala 234:25]
  reg [1:0] states_85_state; // @[elements.scala 234:25]
  reg [1:0] states_86_state; // @[elements.scala 234:25]
  reg [1:0] states_87_state; // @[elements.scala 234:25]
  reg [1:0] states_88_state; // @[elements.scala 234:25]
  reg [1:0] states_89_state; // @[elements.scala 234:25]
  reg [1:0] states_90_state; // @[elements.scala 234:25]
  reg [1:0] states_91_state; // @[elements.scala 234:25]
  reg [1:0] states_92_state; // @[elements.scala 234:25]
  reg [1:0] states_93_state; // @[elements.scala 234:25]
  reg [1:0] states_94_state; // @[elements.scala 234:25]
  reg [1:0] states_95_state; // @[elements.scala 234:25]
  reg [1:0] states_96_state; // @[elements.scala 234:25]
  reg [1:0] states_97_state; // @[elements.scala 234:25]
  reg [1:0] states_98_state; // @[elements.scala 234:25]
  reg [1:0] states_99_state; // @[elements.scala 234:25]
  reg [1:0] states_100_state; // @[elements.scala 234:25]
  reg [1:0] states_101_state; // @[elements.scala 234:25]
  reg [1:0] states_102_state; // @[elements.scala 234:25]
  reg [1:0] states_103_state; // @[elements.scala 234:25]
  reg [1:0] states_104_state; // @[elements.scala 234:25]
  reg [1:0] states_105_state; // @[elements.scala 234:25]
  reg [1:0] states_106_state; // @[elements.scala 234:25]
  reg [1:0] states_107_state; // @[elements.scala 234:25]
  reg [1:0] states_108_state; // @[elements.scala 234:25]
  reg [1:0] states_109_state; // @[elements.scala 234:25]
  reg [1:0] states_110_state; // @[elements.scala 234:25]
  reg [1:0] states_111_state; // @[elements.scala 234:25]
  reg [1:0] states_112_state; // @[elements.scala 234:25]
  reg [1:0] states_113_state; // @[elements.scala 234:25]
  reg [1:0] states_114_state; // @[elements.scala 234:25]
  reg [1:0] states_115_state; // @[elements.scala 234:25]
  reg [1:0] states_116_state; // @[elements.scala 234:25]
  reg [1:0] states_117_state; // @[elements.scala 234:25]
  reg [1:0] states_118_state; // @[elements.scala 234:25]
  reg [1:0] states_119_state; // @[elements.scala 234:25]
  reg [1:0] states_120_state; // @[elements.scala 234:25]
  reg [1:0] states_121_state; // @[elements.scala 234:25]
  reg [1:0] states_122_state; // @[elements.scala 234:25]
  reg [1:0] states_123_state; // @[elements.scala 234:25]
  reg [1:0] states_124_state; // @[elements.scala 234:25]
  reg [1:0] states_125_state; // @[elements.scala 234:25]
  reg [1:0] states_126_state; // @[elements.scala 234:25]
  reg [1:0] states_127_state; // @[elements.scala 234:25]
  reg [1:0] states_128_state; // @[elements.scala 234:25]
  reg [1:0] states_129_state; // @[elements.scala 234:25]
  reg [1:0] states_130_state; // @[elements.scala 234:25]
  reg [1:0] states_131_state; // @[elements.scala 234:25]
  reg [1:0] states_132_state; // @[elements.scala 234:25]
  reg [1:0] states_133_state; // @[elements.scala 234:25]
  reg [1:0] states_134_state; // @[elements.scala 234:25]
  reg [1:0] states_135_state; // @[elements.scala 234:25]
  reg [1:0] states_136_state; // @[elements.scala 234:25]
  reg [1:0] states_137_state; // @[elements.scala 234:25]
  reg [1:0] states_138_state; // @[elements.scala 234:25]
  reg [1:0] states_139_state; // @[elements.scala 234:25]
  reg [1:0] states_140_state; // @[elements.scala 234:25]
  reg [1:0] states_141_state; // @[elements.scala 234:25]
  reg [1:0] states_142_state; // @[elements.scala 234:25]
  reg [1:0] states_143_state; // @[elements.scala 234:25]
  reg [1:0] states_144_state; // @[elements.scala 234:25]
  reg [1:0] states_145_state; // @[elements.scala 234:25]
  reg [1:0] states_146_state; // @[elements.scala 234:25]
  reg [1:0] states_147_state; // @[elements.scala 234:25]
  reg [1:0] states_148_state; // @[elements.scala 234:25]
  reg [1:0] states_149_state; // @[elements.scala 234:25]
  reg [1:0] states_150_state; // @[elements.scala 234:25]
  reg [1:0] states_151_state; // @[elements.scala 234:25]
  reg [1:0] states_152_state; // @[elements.scala 234:25]
  reg [1:0] states_153_state; // @[elements.scala 234:25]
  reg [1:0] states_154_state; // @[elements.scala 234:25]
  reg [1:0] states_155_state; // @[elements.scala 234:25]
  reg [1:0] states_156_state; // @[elements.scala 234:25]
  reg [1:0] states_157_state; // @[elements.scala 234:25]
  reg [1:0] states_158_state; // @[elements.scala 234:25]
  reg [1:0] states_159_state; // @[elements.scala 234:25]
  reg [1:0] states_160_state; // @[elements.scala 234:25]
  reg [1:0] states_161_state; // @[elements.scala 234:25]
  reg [1:0] states_162_state; // @[elements.scala 234:25]
  reg [1:0] states_163_state; // @[elements.scala 234:25]
  reg [1:0] states_164_state; // @[elements.scala 234:25]
  reg [1:0] states_165_state; // @[elements.scala 234:25]
  reg [1:0] states_166_state; // @[elements.scala 234:25]
  reg [1:0] states_167_state; // @[elements.scala 234:25]
  reg [1:0] states_168_state; // @[elements.scala 234:25]
  reg [1:0] states_169_state; // @[elements.scala 234:25]
  reg [1:0] states_170_state; // @[elements.scala 234:25]
  reg [1:0] states_171_state; // @[elements.scala 234:25]
  reg [1:0] states_172_state; // @[elements.scala 234:25]
  reg [1:0] states_173_state; // @[elements.scala 234:25]
  reg [1:0] states_174_state; // @[elements.scala 234:25]
  reg [1:0] states_175_state; // @[elements.scala 234:25]
  reg [1:0] states_176_state; // @[elements.scala 234:25]
  reg [1:0] states_177_state; // @[elements.scala 234:25]
  reg [1:0] states_178_state; // @[elements.scala 234:25]
  reg [1:0] states_179_state; // @[elements.scala 234:25]
  reg [1:0] states_180_state; // @[elements.scala 234:25]
  reg [1:0] states_181_state; // @[elements.scala 234:25]
  reg [1:0] states_182_state; // @[elements.scala 234:25]
  reg [1:0] states_183_state; // @[elements.scala 234:25]
  reg [1:0] states_184_state; // @[elements.scala 234:25]
  reg [1:0] states_185_state; // @[elements.scala 234:25]
  reg [1:0] states_186_state; // @[elements.scala 234:25]
  reg [1:0] states_187_state; // @[elements.scala 234:25]
  reg [1:0] states_188_state; // @[elements.scala 234:25]
  reg [1:0] states_189_state; // @[elements.scala 234:25]
  reg [1:0] states_190_state; // @[elements.scala 234:25]
  reg [1:0] states_191_state; // @[elements.scala 234:25]
  reg [1:0] states_192_state; // @[elements.scala 234:25]
  reg [1:0] states_193_state; // @[elements.scala 234:25]
  reg [1:0] states_194_state; // @[elements.scala 234:25]
  reg [1:0] states_195_state; // @[elements.scala 234:25]
  reg [1:0] states_196_state; // @[elements.scala 234:25]
  reg [1:0] states_197_state; // @[elements.scala 234:25]
  reg [1:0] states_198_state; // @[elements.scala 234:25]
  reg [1:0] states_199_state; // @[elements.scala 234:25]
  reg [1:0] states_200_state; // @[elements.scala 234:25]
  reg [1:0] states_201_state; // @[elements.scala 234:25]
  reg [1:0] states_202_state; // @[elements.scala 234:25]
  reg [1:0] states_203_state; // @[elements.scala 234:25]
  reg [1:0] states_204_state; // @[elements.scala 234:25]
  reg [1:0] states_205_state; // @[elements.scala 234:25]
  reg [1:0] states_206_state; // @[elements.scala 234:25]
  reg [1:0] states_207_state; // @[elements.scala 234:25]
  reg [1:0] states_208_state; // @[elements.scala 234:25]
  reg [1:0] states_209_state; // @[elements.scala 234:25]
  reg [1:0] states_210_state; // @[elements.scala 234:25]
  reg [1:0] states_211_state; // @[elements.scala 234:25]
  reg [1:0] states_212_state; // @[elements.scala 234:25]
  reg [1:0] states_213_state; // @[elements.scala 234:25]
  reg [1:0] states_214_state; // @[elements.scala 234:25]
  reg [1:0] states_215_state; // @[elements.scala 234:25]
  reg [1:0] states_216_state; // @[elements.scala 234:25]
  reg [1:0] states_217_state; // @[elements.scala 234:25]
  reg [1:0] states_218_state; // @[elements.scala 234:25]
  reg [1:0] states_219_state; // @[elements.scala 234:25]
  reg [1:0] states_220_state; // @[elements.scala 234:25]
  reg [1:0] states_221_state; // @[elements.scala 234:25]
  reg [1:0] states_222_state; // @[elements.scala 234:25]
  reg [1:0] states_223_state; // @[elements.scala 234:25]
  reg [1:0] states_224_state; // @[elements.scala 234:25]
  reg [1:0] states_225_state; // @[elements.scala 234:25]
  reg [1:0] states_226_state; // @[elements.scala 234:25]
  reg [1:0] states_227_state; // @[elements.scala 234:25]
  reg [1:0] states_228_state; // @[elements.scala 234:25]
  reg [1:0] states_229_state; // @[elements.scala 234:25]
  reg [1:0] states_230_state; // @[elements.scala 234:25]
  reg [1:0] states_231_state; // @[elements.scala 234:25]
  reg [1:0] states_232_state; // @[elements.scala 234:25]
  reg [1:0] states_233_state; // @[elements.scala 234:25]
  reg [1:0] states_234_state; // @[elements.scala 234:25]
  reg [1:0] states_235_state; // @[elements.scala 234:25]
  reg [1:0] states_236_state; // @[elements.scala 234:25]
  reg [1:0] states_237_state; // @[elements.scala 234:25]
  reg [1:0] states_238_state; // @[elements.scala 234:25]
  reg [1:0] states_239_state; // @[elements.scala 234:25]
  reg [1:0] states_240_state; // @[elements.scala 234:25]
  reg [1:0] states_241_state; // @[elements.scala 234:25]
  reg [1:0] states_242_state; // @[elements.scala 234:25]
  reg [1:0] states_243_state; // @[elements.scala 234:25]
  reg [1:0] states_244_state; // @[elements.scala 234:25]
  reg [1:0] states_245_state; // @[elements.scala 234:25]
  reg [1:0] states_246_state; // @[elements.scala 234:25]
  reg [1:0] states_247_state; // @[elements.scala 234:25]
  reg [1:0] states_248_state; // @[elements.scala 234:25]
  reg [1:0] states_249_state; // @[elements.scala 234:25]
  reg [1:0] states_250_state; // @[elements.scala 234:25]
  reg [1:0] states_251_state; // @[elements.scala 234:25]
  reg [1:0] states_252_state; // @[elements.scala 234:25]
  reg [1:0] states_253_state; // @[elements.scala 234:25]
  reg [1:0] states_254_state; // @[elements.scala 234:25]
  reg [1:0] states_255_state; // @[elements.scala 234:25]
  wire  _T_259 = io_in_1_bits_way != 3'h4; // @[elements.scala 237:91]
  wire  isGet = io_in_1_valid & _T_259; // @[elements.scala 237:66]
  wire  _T_261 = io_in_0_bits_way != 3'h4; // @[elements.scala 243:81]
  wire  isSet_0 = io_in_0_valid & _T_261; // @[elements.scala 243:61]
  wire [8:0] _T_265 = io_in_0_bits_addr[8:3] * 6'h4; // @[elements.scala 244:88]
  wire [8:0] _GEN_768 = {{6'd0}, io_in_0_bits_way}; // @[elements.scala 244:98]
  wire [8:0] _T_267 = _T_265 + _GEN_768; // @[elements.scala 244:98]
  wire [8:0] _T_268 = _T_261 ? _T_267 : 9'h0; // @[elements.scala 244:26]
  wire [7:0] idxSet_0 = _T_268[7:0]; // @[elements.scala 240:23 elements.scala 244:20]
  wire [8:0] _T_271 = io_in_1_bits_addr[8:3] * 6'h4; // @[elements.scala 253:91]
  wire [8:0] _GEN_769 = {{6'd0}, io_in_1_bits_way}; // @[elements.scala 253:101]
  wire [8:0] _T_273 = _T_271 + _GEN_769; // @[elements.scala 253:101]
  wire [8:0] _T_274 = _T_259 ? _T_273 : 9'h0; // @[elements.scala 253:19]
  wire [7:0] idxGet = _T_274[7:0]; // @[elements.scala 239:22 elements.scala 253:12]
  wire [1:0] _GEN_513 = 8'h1 == idxGet ? states_1_state : states_0_state; // @[elements.scala 254:17]
  wire [1:0] _GEN_514 = 8'h2 == idxGet ? states_2_state : _GEN_513; // @[elements.scala 254:17]
  wire [1:0] _GEN_515 = 8'h3 == idxGet ? states_3_state : _GEN_514; // @[elements.scala 254:17]
  wire [1:0] _GEN_516 = 8'h4 == idxGet ? states_4_state : _GEN_515; // @[elements.scala 254:17]
  wire [1:0] _GEN_517 = 8'h5 == idxGet ? states_5_state : _GEN_516; // @[elements.scala 254:17]
  wire [1:0] _GEN_518 = 8'h6 == idxGet ? states_6_state : _GEN_517; // @[elements.scala 254:17]
  wire [1:0] _GEN_519 = 8'h7 == idxGet ? states_7_state : _GEN_518; // @[elements.scala 254:17]
  wire [1:0] _GEN_520 = 8'h8 == idxGet ? states_8_state : _GEN_519; // @[elements.scala 254:17]
  wire [1:0] _GEN_521 = 8'h9 == idxGet ? states_9_state : _GEN_520; // @[elements.scala 254:17]
  wire [1:0] _GEN_522 = 8'ha == idxGet ? states_10_state : _GEN_521; // @[elements.scala 254:17]
  wire [1:0] _GEN_523 = 8'hb == idxGet ? states_11_state : _GEN_522; // @[elements.scala 254:17]
  wire [1:0] _GEN_524 = 8'hc == idxGet ? states_12_state : _GEN_523; // @[elements.scala 254:17]
  wire [1:0] _GEN_525 = 8'hd == idxGet ? states_13_state : _GEN_524; // @[elements.scala 254:17]
  wire [1:0] _GEN_526 = 8'he == idxGet ? states_14_state : _GEN_525; // @[elements.scala 254:17]
  wire [1:0] _GEN_527 = 8'hf == idxGet ? states_15_state : _GEN_526; // @[elements.scala 254:17]
  wire [1:0] _GEN_528 = 8'h10 == idxGet ? states_16_state : _GEN_527; // @[elements.scala 254:17]
  wire [1:0] _GEN_529 = 8'h11 == idxGet ? states_17_state : _GEN_528; // @[elements.scala 254:17]
  wire [1:0] _GEN_530 = 8'h12 == idxGet ? states_18_state : _GEN_529; // @[elements.scala 254:17]
  wire [1:0] _GEN_531 = 8'h13 == idxGet ? states_19_state : _GEN_530; // @[elements.scala 254:17]
  wire [1:0] _GEN_532 = 8'h14 == idxGet ? states_20_state : _GEN_531; // @[elements.scala 254:17]
  wire [1:0] _GEN_533 = 8'h15 == idxGet ? states_21_state : _GEN_532; // @[elements.scala 254:17]
  wire [1:0] _GEN_534 = 8'h16 == idxGet ? states_22_state : _GEN_533; // @[elements.scala 254:17]
  wire [1:0] _GEN_535 = 8'h17 == idxGet ? states_23_state : _GEN_534; // @[elements.scala 254:17]
  wire [1:0] _GEN_536 = 8'h18 == idxGet ? states_24_state : _GEN_535; // @[elements.scala 254:17]
  wire [1:0] _GEN_537 = 8'h19 == idxGet ? states_25_state : _GEN_536; // @[elements.scala 254:17]
  wire [1:0] _GEN_538 = 8'h1a == idxGet ? states_26_state : _GEN_537; // @[elements.scala 254:17]
  wire [1:0] _GEN_539 = 8'h1b == idxGet ? states_27_state : _GEN_538; // @[elements.scala 254:17]
  wire [1:0] _GEN_540 = 8'h1c == idxGet ? states_28_state : _GEN_539; // @[elements.scala 254:17]
  wire [1:0] _GEN_541 = 8'h1d == idxGet ? states_29_state : _GEN_540; // @[elements.scala 254:17]
  wire [1:0] _GEN_542 = 8'h1e == idxGet ? states_30_state : _GEN_541; // @[elements.scala 254:17]
  wire [1:0] _GEN_543 = 8'h1f == idxGet ? states_31_state : _GEN_542; // @[elements.scala 254:17]
  wire [1:0] _GEN_544 = 8'h20 == idxGet ? states_32_state : _GEN_543; // @[elements.scala 254:17]
  wire [1:0] _GEN_545 = 8'h21 == idxGet ? states_33_state : _GEN_544; // @[elements.scala 254:17]
  wire [1:0] _GEN_546 = 8'h22 == idxGet ? states_34_state : _GEN_545; // @[elements.scala 254:17]
  wire [1:0] _GEN_547 = 8'h23 == idxGet ? states_35_state : _GEN_546; // @[elements.scala 254:17]
  wire [1:0] _GEN_548 = 8'h24 == idxGet ? states_36_state : _GEN_547; // @[elements.scala 254:17]
  wire [1:0] _GEN_549 = 8'h25 == idxGet ? states_37_state : _GEN_548; // @[elements.scala 254:17]
  wire [1:0] _GEN_550 = 8'h26 == idxGet ? states_38_state : _GEN_549; // @[elements.scala 254:17]
  wire [1:0] _GEN_551 = 8'h27 == idxGet ? states_39_state : _GEN_550; // @[elements.scala 254:17]
  wire [1:0] _GEN_552 = 8'h28 == idxGet ? states_40_state : _GEN_551; // @[elements.scala 254:17]
  wire [1:0] _GEN_553 = 8'h29 == idxGet ? states_41_state : _GEN_552; // @[elements.scala 254:17]
  wire [1:0] _GEN_554 = 8'h2a == idxGet ? states_42_state : _GEN_553; // @[elements.scala 254:17]
  wire [1:0] _GEN_555 = 8'h2b == idxGet ? states_43_state : _GEN_554; // @[elements.scala 254:17]
  wire [1:0] _GEN_556 = 8'h2c == idxGet ? states_44_state : _GEN_555; // @[elements.scala 254:17]
  wire [1:0] _GEN_557 = 8'h2d == idxGet ? states_45_state : _GEN_556; // @[elements.scala 254:17]
  wire [1:0] _GEN_558 = 8'h2e == idxGet ? states_46_state : _GEN_557; // @[elements.scala 254:17]
  wire [1:0] _GEN_559 = 8'h2f == idxGet ? states_47_state : _GEN_558; // @[elements.scala 254:17]
  wire [1:0] _GEN_560 = 8'h30 == idxGet ? states_48_state : _GEN_559; // @[elements.scala 254:17]
  wire [1:0] _GEN_561 = 8'h31 == idxGet ? states_49_state : _GEN_560; // @[elements.scala 254:17]
  wire [1:0] _GEN_562 = 8'h32 == idxGet ? states_50_state : _GEN_561; // @[elements.scala 254:17]
  wire [1:0] _GEN_563 = 8'h33 == idxGet ? states_51_state : _GEN_562; // @[elements.scala 254:17]
  wire [1:0] _GEN_564 = 8'h34 == idxGet ? states_52_state : _GEN_563; // @[elements.scala 254:17]
  wire [1:0] _GEN_565 = 8'h35 == idxGet ? states_53_state : _GEN_564; // @[elements.scala 254:17]
  wire [1:0] _GEN_566 = 8'h36 == idxGet ? states_54_state : _GEN_565; // @[elements.scala 254:17]
  wire [1:0] _GEN_567 = 8'h37 == idxGet ? states_55_state : _GEN_566; // @[elements.scala 254:17]
  wire [1:0] _GEN_568 = 8'h38 == idxGet ? states_56_state : _GEN_567; // @[elements.scala 254:17]
  wire [1:0] _GEN_569 = 8'h39 == idxGet ? states_57_state : _GEN_568; // @[elements.scala 254:17]
  wire [1:0] _GEN_570 = 8'h3a == idxGet ? states_58_state : _GEN_569; // @[elements.scala 254:17]
  wire [1:0] _GEN_571 = 8'h3b == idxGet ? states_59_state : _GEN_570; // @[elements.scala 254:17]
  wire [1:0] _GEN_572 = 8'h3c == idxGet ? states_60_state : _GEN_571; // @[elements.scala 254:17]
  wire [1:0] _GEN_573 = 8'h3d == idxGet ? states_61_state : _GEN_572; // @[elements.scala 254:17]
  wire [1:0] _GEN_574 = 8'h3e == idxGet ? states_62_state : _GEN_573; // @[elements.scala 254:17]
  wire [1:0] _GEN_575 = 8'h3f == idxGet ? states_63_state : _GEN_574; // @[elements.scala 254:17]
  wire [1:0] _GEN_576 = 8'h40 == idxGet ? states_64_state : _GEN_575; // @[elements.scala 254:17]
  wire [1:0] _GEN_577 = 8'h41 == idxGet ? states_65_state : _GEN_576; // @[elements.scala 254:17]
  wire [1:0] _GEN_578 = 8'h42 == idxGet ? states_66_state : _GEN_577; // @[elements.scala 254:17]
  wire [1:0] _GEN_579 = 8'h43 == idxGet ? states_67_state : _GEN_578; // @[elements.scala 254:17]
  wire [1:0] _GEN_580 = 8'h44 == idxGet ? states_68_state : _GEN_579; // @[elements.scala 254:17]
  wire [1:0] _GEN_581 = 8'h45 == idxGet ? states_69_state : _GEN_580; // @[elements.scala 254:17]
  wire [1:0] _GEN_582 = 8'h46 == idxGet ? states_70_state : _GEN_581; // @[elements.scala 254:17]
  wire [1:0] _GEN_583 = 8'h47 == idxGet ? states_71_state : _GEN_582; // @[elements.scala 254:17]
  wire [1:0] _GEN_584 = 8'h48 == idxGet ? states_72_state : _GEN_583; // @[elements.scala 254:17]
  wire [1:0] _GEN_585 = 8'h49 == idxGet ? states_73_state : _GEN_584; // @[elements.scala 254:17]
  wire [1:0] _GEN_586 = 8'h4a == idxGet ? states_74_state : _GEN_585; // @[elements.scala 254:17]
  wire [1:0] _GEN_587 = 8'h4b == idxGet ? states_75_state : _GEN_586; // @[elements.scala 254:17]
  wire [1:0] _GEN_588 = 8'h4c == idxGet ? states_76_state : _GEN_587; // @[elements.scala 254:17]
  wire [1:0] _GEN_589 = 8'h4d == idxGet ? states_77_state : _GEN_588; // @[elements.scala 254:17]
  wire [1:0] _GEN_590 = 8'h4e == idxGet ? states_78_state : _GEN_589; // @[elements.scala 254:17]
  wire [1:0] _GEN_591 = 8'h4f == idxGet ? states_79_state : _GEN_590; // @[elements.scala 254:17]
  wire [1:0] _GEN_592 = 8'h50 == idxGet ? states_80_state : _GEN_591; // @[elements.scala 254:17]
  wire [1:0] _GEN_593 = 8'h51 == idxGet ? states_81_state : _GEN_592; // @[elements.scala 254:17]
  wire [1:0] _GEN_594 = 8'h52 == idxGet ? states_82_state : _GEN_593; // @[elements.scala 254:17]
  wire [1:0] _GEN_595 = 8'h53 == idxGet ? states_83_state : _GEN_594; // @[elements.scala 254:17]
  wire [1:0] _GEN_596 = 8'h54 == idxGet ? states_84_state : _GEN_595; // @[elements.scala 254:17]
  wire [1:0] _GEN_597 = 8'h55 == idxGet ? states_85_state : _GEN_596; // @[elements.scala 254:17]
  wire [1:0] _GEN_598 = 8'h56 == idxGet ? states_86_state : _GEN_597; // @[elements.scala 254:17]
  wire [1:0] _GEN_599 = 8'h57 == idxGet ? states_87_state : _GEN_598; // @[elements.scala 254:17]
  wire [1:0] _GEN_600 = 8'h58 == idxGet ? states_88_state : _GEN_599; // @[elements.scala 254:17]
  wire [1:0] _GEN_601 = 8'h59 == idxGet ? states_89_state : _GEN_600; // @[elements.scala 254:17]
  wire [1:0] _GEN_602 = 8'h5a == idxGet ? states_90_state : _GEN_601; // @[elements.scala 254:17]
  wire [1:0] _GEN_603 = 8'h5b == idxGet ? states_91_state : _GEN_602; // @[elements.scala 254:17]
  wire [1:0] _GEN_604 = 8'h5c == idxGet ? states_92_state : _GEN_603; // @[elements.scala 254:17]
  wire [1:0] _GEN_605 = 8'h5d == idxGet ? states_93_state : _GEN_604; // @[elements.scala 254:17]
  wire [1:0] _GEN_606 = 8'h5e == idxGet ? states_94_state : _GEN_605; // @[elements.scala 254:17]
  wire [1:0] _GEN_607 = 8'h5f == idxGet ? states_95_state : _GEN_606; // @[elements.scala 254:17]
  wire [1:0] _GEN_608 = 8'h60 == idxGet ? states_96_state : _GEN_607; // @[elements.scala 254:17]
  wire [1:0] _GEN_609 = 8'h61 == idxGet ? states_97_state : _GEN_608; // @[elements.scala 254:17]
  wire [1:0] _GEN_610 = 8'h62 == idxGet ? states_98_state : _GEN_609; // @[elements.scala 254:17]
  wire [1:0] _GEN_611 = 8'h63 == idxGet ? states_99_state : _GEN_610; // @[elements.scala 254:17]
  wire [1:0] _GEN_612 = 8'h64 == idxGet ? states_100_state : _GEN_611; // @[elements.scala 254:17]
  wire [1:0] _GEN_613 = 8'h65 == idxGet ? states_101_state : _GEN_612; // @[elements.scala 254:17]
  wire [1:0] _GEN_614 = 8'h66 == idxGet ? states_102_state : _GEN_613; // @[elements.scala 254:17]
  wire [1:0] _GEN_615 = 8'h67 == idxGet ? states_103_state : _GEN_614; // @[elements.scala 254:17]
  wire [1:0] _GEN_616 = 8'h68 == idxGet ? states_104_state : _GEN_615; // @[elements.scala 254:17]
  wire [1:0] _GEN_617 = 8'h69 == idxGet ? states_105_state : _GEN_616; // @[elements.scala 254:17]
  wire [1:0] _GEN_618 = 8'h6a == idxGet ? states_106_state : _GEN_617; // @[elements.scala 254:17]
  wire [1:0] _GEN_619 = 8'h6b == idxGet ? states_107_state : _GEN_618; // @[elements.scala 254:17]
  wire [1:0] _GEN_620 = 8'h6c == idxGet ? states_108_state : _GEN_619; // @[elements.scala 254:17]
  wire [1:0] _GEN_621 = 8'h6d == idxGet ? states_109_state : _GEN_620; // @[elements.scala 254:17]
  wire [1:0] _GEN_622 = 8'h6e == idxGet ? states_110_state : _GEN_621; // @[elements.scala 254:17]
  wire [1:0] _GEN_623 = 8'h6f == idxGet ? states_111_state : _GEN_622; // @[elements.scala 254:17]
  wire [1:0] _GEN_624 = 8'h70 == idxGet ? states_112_state : _GEN_623; // @[elements.scala 254:17]
  wire [1:0] _GEN_625 = 8'h71 == idxGet ? states_113_state : _GEN_624; // @[elements.scala 254:17]
  wire [1:0] _GEN_626 = 8'h72 == idxGet ? states_114_state : _GEN_625; // @[elements.scala 254:17]
  wire [1:0] _GEN_627 = 8'h73 == idxGet ? states_115_state : _GEN_626; // @[elements.scala 254:17]
  wire [1:0] _GEN_628 = 8'h74 == idxGet ? states_116_state : _GEN_627; // @[elements.scala 254:17]
  wire [1:0] _GEN_629 = 8'h75 == idxGet ? states_117_state : _GEN_628; // @[elements.scala 254:17]
  wire [1:0] _GEN_630 = 8'h76 == idxGet ? states_118_state : _GEN_629; // @[elements.scala 254:17]
  wire [1:0] _GEN_631 = 8'h77 == idxGet ? states_119_state : _GEN_630; // @[elements.scala 254:17]
  wire [1:0] _GEN_632 = 8'h78 == idxGet ? states_120_state : _GEN_631; // @[elements.scala 254:17]
  wire [1:0] _GEN_633 = 8'h79 == idxGet ? states_121_state : _GEN_632; // @[elements.scala 254:17]
  wire [1:0] _GEN_634 = 8'h7a == idxGet ? states_122_state : _GEN_633; // @[elements.scala 254:17]
  wire [1:0] _GEN_635 = 8'h7b == idxGet ? states_123_state : _GEN_634; // @[elements.scala 254:17]
  wire [1:0] _GEN_636 = 8'h7c == idxGet ? states_124_state : _GEN_635; // @[elements.scala 254:17]
  wire [1:0] _GEN_637 = 8'h7d == idxGet ? states_125_state : _GEN_636; // @[elements.scala 254:17]
  wire [1:0] _GEN_638 = 8'h7e == idxGet ? states_126_state : _GEN_637; // @[elements.scala 254:17]
  wire [1:0] _GEN_639 = 8'h7f == idxGet ? states_127_state : _GEN_638; // @[elements.scala 254:17]
  wire [1:0] _GEN_640 = 8'h80 == idxGet ? states_128_state : _GEN_639; // @[elements.scala 254:17]
  wire [1:0] _GEN_641 = 8'h81 == idxGet ? states_129_state : _GEN_640; // @[elements.scala 254:17]
  wire [1:0] _GEN_642 = 8'h82 == idxGet ? states_130_state : _GEN_641; // @[elements.scala 254:17]
  wire [1:0] _GEN_643 = 8'h83 == idxGet ? states_131_state : _GEN_642; // @[elements.scala 254:17]
  wire [1:0] _GEN_644 = 8'h84 == idxGet ? states_132_state : _GEN_643; // @[elements.scala 254:17]
  wire [1:0] _GEN_645 = 8'h85 == idxGet ? states_133_state : _GEN_644; // @[elements.scala 254:17]
  wire [1:0] _GEN_646 = 8'h86 == idxGet ? states_134_state : _GEN_645; // @[elements.scala 254:17]
  wire [1:0] _GEN_647 = 8'h87 == idxGet ? states_135_state : _GEN_646; // @[elements.scala 254:17]
  wire [1:0] _GEN_648 = 8'h88 == idxGet ? states_136_state : _GEN_647; // @[elements.scala 254:17]
  wire [1:0] _GEN_649 = 8'h89 == idxGet ? states_137_state : _GEN_648; // @[elements.scala 254:17]
  wire [1:0] _GEN_650 = 8'h8a == idxGet ? states_138_state : _GEN_649; // @[elements.scala 254:17]
  wire [1:0] _GEN_651 = 8'h8b == idxGet ? states_139_state : _GEN_650; // @[elements.scala 254:17]
  wire [1:0] _GEN_652 = 8'h8c == idxGet ? states_140_state : _GEN_651; // @[elements.scala 254:17]
  wire [1:0] _GEN_653 = 8'h8d == idxGet ? states_141_state : _GEN_652; // @[elements.scala 254:17]
  wire [1:0] _GEN_654 = 8'h8e == idxGet ? states_142_state : _GEN_653; // @[elements.scala 254:17]
  wire [1:0] _GEN_655 = 8'h8f == idxGet ? states_143_state : _GEN_654; // @[elements.scala 254:17]
  wire [1:0] _GEN_656 = 8'h90 == idxGet ? states_144_state : _GEN_655; // @[elements.scala 254:17]
  wire [1:0] _GEN_657 = 8'h91 == idxGet ? states_145_state : _GEN_656; // @[elements.scala 254:17]
  wire [1:0] _GEN_658 = 8'h92 == idxGet ? states_146_state : _GEN_657; // @[elements.scala 254:17]
  wire [1:0] _GEN_659 = 8'h93 == idxGet ? states_147_state : _GEN_658; // @[elements.scala 254:17]
  wire [1:0] _GEN_660 = 8'h94 == idxGet ? states_148_state : _GEN_659; // @[elements.scala 254:17]
  wire [1:0] _GEN_661 = 8'h95 == idxGet ? states_149_state : _GEN_660; // @[elements.scala 254:17]
  wire [1:0] _GEN_662 = 8'h96 == idxGet ? states_150_state : _GEN_661; // @[elements.scala 254:17]
  wire [1:0] _GEN_663 = 8'h97 == idxGet ? states_151_state : _GEN_662; // @[elements.scala 254:17]
  wire [1:0] _GEN_664 = 8'h98 == idxGet ? states_152_state : _GEN_663; // @[elements.scala 254:17]
  wire [1:0] _GEN_665 = 8'h99 == idxGet ? states_153_state : _GEN_664; // @[elements.scala 254:17]
  wire [1:0] _GEN_666 = 8'h9a == idxGet ? states_154_state : _GEN_665; // @[elements.scala 254:17]
  wire [1:0] _GEN_667 = 8'h9b == idxGet ? states_155_state : _GEN_666; // @[elements.scala 254:17]
  wire [1:0] _GEN_668 = 8'h9c == idxGet ? states_156_state : _GEN_667; // @[elements.scala 254:17]
  wire [1:0] _GEN_669 = 8'h9d == idxGet ? states_157_state : _GEN_668; // @[elements.scala 254:17]
  wire [1:0] _GEN_670 = 8'h9e == idxGet ? states_158_state : _GEN_669; // @[elements.scala 254:17]
  wire [1:0] _GEN_671 = 8'h9f == idxGet ? states_159_state : _GEN_670; // @[elements.scala 254:17]
  wire [1:0] _GEN_672 = 8'ha0 == idxGet ? states_160_state : _GEN_671; // @[elements.scala 254:17]
  wire [1:0] _GEN_673 = 8'ha1 == idxGet ? states_161_state : _GEN_672; // @[elements.scala 254:17]
  wire [1:0] _GEN_674 = 8'ha2 == idxGet ? states_162_state : _GEN_673; // @[elements.scala 254:17]
  wire [1:0] _GEN_675 = 8'ha3 == idxGet ? states_163_state : _GEN_674; // @[elements.scala 254:17]
  wire [1:0] _GEN_676 = 8'ha4 == idxGet ? states_164_state : _GEN_675; // @[elements.scala 254:17]
  wire [1:0] _GEN_677 = 8'ha5 == idxGet ? states_165_state : _GEN_676; // @[elements.scala 254:17]
  wire [1:0] _GEN_678 = 8'ha6 == idxGet ? states_166_state : _GEN_677; // @[elements.scala 254:17]
  wire [1:0] _GEN_679 = 8'ha7 == idxGet ? states_167_state : _GEN_678; // @[elements.scala 254:17]
  wire [1:0] _GEN_680 = 8'ha8 == idxGet ? states_168_state : _GEN_679; // @[elements.scala 254:17]
  wire [1:0] _GEN_681 = 8'ha9 == idxGet ? states_169_state : _GEN_680; // @[elements.scala 254:17]
  wire [1:0] _GEN_682 = 8'haa == idxGet ? states_170_state : _GEN_681; // @[elements.scala 254:17]
  wire [1:0] _GEN_683 = 8'hab == idxGet ? states_171_state : _GEN_682; // @[elements.scala 254:17]
  wire [1:0] _GEN_684 = 8'hac == idxGet ? states_172_state : _GEN_683; // @[elements.scala 254:17]
  wire [1:0] _GEN_685 = 8'had == idxGet ? states_173_state : _GEN_684; // @[elements.scala 254:17]
  wire [1:0] _GEN_686 = 8'hae == idxGet ? states_174_state : _GEN_685; // @[elements.scala 254:17]
  wire [1:0] _GEN_687 = 8'haf == idxGet ? states_175_state : _GEN_686; // @[elements.scala 254:17]
  wire [1:0] _GEN_688 = 8'hb0 == idxGet ? states_176_state : _GEN_687; // @[elements.scala 254:17]
  wire [1:0] _GEN_689 = 8'hb1 == idxGet ? states_177_state : _GEN_688; // @[elements.scala 254:17]
  wire [1:0] _GEN_690 = 8'hb2 == idxGet ? states_178_state : _GEN_689; // @[elements.scala 254:17]
  wire [1:0] _GEN_691 = 8'hb3 == idxGet ? states_179_state : _GEN_690; // @[elements.scala 254:17]
  wire [1:0] _GEN_692 = 8'hb4 == idxGet ? states_180_state : _GEN_691; // @[elements.scala 254:17]
  wire [1:0] _GEN_693 = 8'hb5 == idxGet ? states_181_state : _GEN_692; // @[elements.scala 254:17]
  wire [1:0] _GEN_694 = 8'hb6 == idxGet ? states_182_state : _GEN_693; // @[elements.scala 254:17]
  wire [1:0] _GEN_695 = 8'hb7 == idxGet ? states_183_state : _GEN_694; // @[elements.scala 254:17]
  wire [1:0] _GEN_696 = 8'hb8 == idxGet ? states_184_state : _GEN_695; // @[elements.scala 254:17]
  wire [1:0] _GEN_697 = 8'hb9 == idxGet ? states_185_state : _GEN_696; // @[elements.scala 254:17]
  wire [1:0] _GEN_698 = 8'hba == idxGet ? states_186_state : _GEN_697; // @[elements.scala 254:17]
  wire [1:0] _GEN_699 = 8'hbb == idxGet ? states_187_state : _GEN_698; // @[elements.scala 254:17]
  wire [1:0] _GEN_700 = 8'hbc == idxGet ? states_188_state : _GEN_699; // @[elements.scala 254:17]
  wire [1:0] _GEN_701 = 8'hbd == idxGet ? states_189_state : _GEN_700; // @[elements.scala 254:17]
  wire [1:0] _GEN_702 = 8'hbe == idxGet ? states_190_state : _GEN_701; // @[elements.scala 254:17]
  wire [1:0] _GEN_703 = 8'hbf == idxGet ? states_191_state : _GEN_702; // @[elements.scala 254:17]
  wire [1:0] _GEN_704 = 8'hc0 == idxGet ? states_192_state : _GEN_703; // @[elements.scala 254:17]
  wire [1:0] _GEN_705 = 8'hc1 == idxGet ? states_193_state : _GEN_704; // @[elements.scala 254:17]
  wire [1:0] _GEN_706 = 8'hc2 == idxGet ? states_194_state : _GEN_705; // @[elements.scala 254:17]
  wire [1:0] _GEN_707 = 8'hc3 == idxGet ? states_195_state : _GEN_706; // @[elements.scala 254:17]
  wire [1:0] _GEN_708 = 8'hc4 == idxGet ? states_196_state : _GEN_707; // @[elements.scala 254:17]
  wire [1:0] _GEN_709 = 8'hc5 == idxGet ? states_197_state : _GEN_708; // @[elements.scala 254:17]
  wire [1:0] _GEN_710 = 8'hc6 == idxGet ? states_198_state : _GEN_709; // @[elements.scala 254:17]
  wire [1:0] _GEN_711 = 8'hc7 == idxGet ? states_199_state : _GEN_710; // @[elements.scala 254:17]
  wire [1:0] _GEN_712 = 8'hc8 == idxGet ? states_200_state : _GEN_711; // @[elements.scala 254:17]
  wire [1:0] _GEN_713 = 8'hc9 == idxGet ? states_201_state : _GEN_712; // @[elements.scala 254:17]
  wire [1:0] _GEN_714 = 8'hca == idxGet ? states_202_state : _GEN_713; // @[elements.scala 254:17]
  wire [1:0] _GEN_715 = 8'hcb == idxGet ? states_203_state : _GEN_714; // @[elements.scala 254:17]
  wire [1:0] _GEN_716 = 8'hcc == idxGet ? states_204_state : _GEN_715; // @[elements.scala 254:17]
  wire [1:0] _GEN_717 = 8'hcd == idxGet ? states_205_state : _GEN_716; // @[elements.scala 254:17]
  wire [1:0] _GEN_718 = 8'hce == idxGet ? states_206_state : _GEN_717; // @[elements.scala 254:17]
  wire [1:0] _GEN_719 = 8'hcf == idxGet ? states_207_state : _GEN_718; // @[elements.scala 254:17]
  wire [1:0] _GEN_720 = 8'hd0 == idxGet ? states_208_state : _GEN_719; // @[elements.scala 254:17]
  wire [1:0] _GEN_721 = 8'hd1 == idxGet ? states_209_state : _GEN_720; // @[elements.scala 254:17]
  wire [1:0] _GEN_722 = 8'hd2 == idxGet ? states_210_state : _GEN_721; // @[elements.scala 254:17]
  wire [1:0] _GEN_723 = 8'hd3 == idxGet ? states_211_state : _GEN_722; // @[elements.scala 254:17]
  wire [1:0] _GEN_724 = 8'hd4 == idxGet ? states_212_state : _GEN_723; // @[elements.scala 254:17]
  wire [1:0] _GEN_725 = 8'hd5 == idxGet ? states_213_state : _GEN_724; // @[elements.scala 254:17]
  wire [1:0] _GEN_726 = 8'hd6 == idxGet ? states_214_state : _GEN_725; // @[elements.scala 254:17]
  wire [1:0] _GEN_727 = 8'hd7 == idxGet ? states_215_state : _GEN_726; // @[elements.scala 254:17]
  wire [1:0] _GEN_728 = 8'hd8 == idxGet ? states_216_state : _GEN_727; // @[elements.scala 254:17]
  wire [1:0] _GEN_729 = 8'hd9 == idxGet ? states_217_state : _GEN_728; // @[elements.scala 254:17]
  wire [1:0] _GEN_730 = 8'hda == idxGet ? states_218_state : _GEN_729; // @[elements.scala 254:17]
  wire [1:0] _GEN_731 = 8'hdb == idxGet ? states_219_state : _GEN_730; // @[elements.scala 254:17]
  wire [1:0] _GEN_732 = 8'hdc == idxGet ? states_220_state : _GEN_731; // @[elements.scala 254:17]
  wire [1:0] _GEN_733 = 8'hdd == idxGet ? states_221_state : _GEN_732; // @[elements.scala 254:17]
  wire [1:0] _GEN_734 = 8'hde == idxGet ? states_222_state : _GEN_733; // @[elements.scala 254:17]
  wire [1:0] _GEN_735 = 8'hdf == idxGet ? states_223_state : _GEN_734; // @[elements.scala 254:17]
  wire [1:0] _GEN_736 = 8'he0 == idxGet ? states_224_state : _GEN_735; // @[elements.scala 254:17]
  wire [1:0] _GEN_737 = 8'he1 == idxGet ? states_225_state : _GEN_736; // @[elements.scala 254:17]
  wire [1:0] _GEN_738 = 8'he2 == idxGet ? states_226_state : _GEN_737; // @[elements.scala 254:17]
  wire [1:0] _GEN_739 = 8'he3 == idxGet ? states_227_state : _GEN_738; // @[elements.scala 254:17]
  wire [1:0] _GEN_740 = 8'he4 == idxGet ? states_228_state : _GEN_739; // @[elements.scala 254:17]
  wire [1:0] _GEN_741 = 8'he5 == idxGet ? states_229_state : _GEN_740; // @[elements.scala 254:17]
  wire [1:0] _GEN_742 = 8'he6 == idxGet ? states_230_state : _GEN_741; // @[elements.scala 254:17]
  wire [1:0] _GEN_743 = 8'he7 == idxGet ? states_231_state : _GEN_742; // @[elements.scala 254:17]
  wire [1:0] _GEN_744 = 8'he8 == idxGet ? states_232_state : _GEN_743; // @[elements.scala 254:17]
  wire [1:0] _GEN_745 = 8'he9 == idxGet ? states_233_state : _GEN_744; // @[elements.scala 254:17]
  wire [1:0] _GEN_746 = 8'hea == idxGet ? states_234_state : _GEN_745; // @[elements.scala 254:17]
  wire [1:0] _GEN_747 = 8'heb == idxGet ? states_235_state : _GEN_746; // @[elements.scala 254:17]
  wire [1:0] _GEN_748 = 8'hec == idxGet ? states_236_state : _GEN_747; // @[elements.scala 254:17]
  wire [1:0] _GEN_749 = 8'hed == idxGet ? states_237_state : _GEN_748; // @[elements.scala 254:17]
  wire [1:0] _GEN_750 = 8'hee == idxGet ? states_238_state : _GEN_749; // @[elements.scala 254:17]
  wire [1:0] _GEN_751 = 8'hef == idxGet ? states_239_state : _GEN_750; // @[elements.scala 254:17]
  wire [1:0] _GEN_752 = 8'hf0 == idxGet ? states_240_state : _GEN_751; // @[elements.scala 254:17]
  wire [1:0] _GEN_753 = 8'hf1 == idxGet ? states_241_state : _GEN_752; // @[elements.scala 254:17]
  wire [1:0] _GEN_754 = 8'hf2 == idxGet ? states_242_state : _GEN_753; // @[elements.scala 254:17]
  wire [1:0] _GEN_755 = 8'hf3 == idxGet ? states_243_state : _GEN_754; // @[elements.scala 254:17]
  wire [1:0] _GEN_756 = 8'hf4 == idxGet ? states_244_state : _GEN_755; // @[elements.scala 254:17]
  wire [1:0] _GEN_757 = 8'hf5 == idxGet ? states_245_state : _GEN_756; // @[elements.scala 254:17]
  wire [1:0] _GEN_758 = 8'hf6 == idxGet ? states_246_state : _GEN_757; // @[elements.scala 254:17]
  wire [1:0] _GEN_759 = 8'hf7 == idxGet ? states_247_state : _GEN_758; // @[elements.scala 254:17]
  wire [1:0] _GEN_760 = 8'hf8 == idxGet ? states_248_state : _GEN_759; // @[elements.scala 254:17]
  wire [1:0] _GEN_761 = 8'hf9 == idxGet ? states_249_state : _GEN_760; // @[elements.scala 254:17]
  wire [1:0] _GEN_762 = 8'hfa == idxGet ? states_250_state : _GEN_761; // @[elements.scala 254:17]
  wire [1:0] _GEN_763 = 8'hfb == idxGet ? states_251_state : _GEN_762; // @[elements.scala 254:17]
  wire [1:0] _GEN_764 = 8'hfc == idxGet ? states_252_state : _GEN_763; // @[elements.scala 254:17]
  wire [1:0] _GEN_765 = 8'hfd == idxGet ? states_253_state : _GEN_764; // @[elements.scala 254:17]
  wire [1:0] _GEN_766 = 8'hfe == idxGet ? states_254_state : _GEN_765; // @[elements.scala 254:17]
  assign io_out_valid = _T_259 & isGet; // @[elements.scala 255:18]
  assign io_out_bits_state = 8'hff == idxGet ? states_255_state : _GEN_766; // @[elements.scala 254:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  states_0_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  states_1_state = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  states_2_state = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  states_3_state = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  states_4_state = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  states_5_state = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  states_6_state = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  states_7_state = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  states_8_state = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  states_9_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  states_10_state = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  states_11_state = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  states_12_state = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  states_13_state = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  states_14_state = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  states_15_state = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  states_16_state = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  states_17_state = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  states_18_state = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  states_19_state = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  states_20_state = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  states_21_state = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  states_22_state = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  states_23_state = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  states_24_state = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  states_25_state = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  states_26_state = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  states_27_state = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  states_28_state = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  states_29_state = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  states_30_state = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  states_31_state = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  states_32_state = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  states_33_state = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  states_34_state = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  states_35_state = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  states_36_state = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  states_37_state = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  states_38_state = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  states_39_state = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  states_40_state = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  states_41_state = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  states_42_state = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  states_43_state = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  states_44_state = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  states_45_state = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  states_46_state = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  states_47_state = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  states_48_state = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  states_49_state = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  states_50_state = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  states_51_state = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  states_52_state = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  states_53_state = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  states_54_state = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  states_55_state = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  states_56_state = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  states_57_state = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  states_58_state = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  states_59_state = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  states_60_state = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  states_61_state = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  states_62_state = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  states_63_state = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  states_64_state = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  states_65_state = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  states_66_state = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  states_67_state = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  states_68_state = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  states_69_state = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  states_70_state = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  states_71_state = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  states_72_state = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  states_73_state = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  states_74_state = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  states_75_state = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  states_76_state = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  states_77_state = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  states_78_state = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  states_79_state = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  states_80_state = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  states_81_state = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  states_82_state = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  states_83_state = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  states_84_state = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  states_85_state = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  states_86_state = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  states_87_state = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  states_88_state = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  states_89_state = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  states_90_state = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  states_91_state = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  states_92_state = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  states_93_state = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  states_94_state = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  states_95_state = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  states_96_state = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  states_97_state = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  states_98_state = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  states_99_state = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  states_100_state = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  states_101_state = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  states_102_state = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  states_103_state = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  states_104_state = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  states_105_state = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  states_106_state = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  states_107_state = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  states_108_state = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  states_109_state = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  states_110_state = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  states_111_state = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  states_112_state = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  states_113_state = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  states_114_state = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  states_115_state = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  states_116_state = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  states_117_state = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  states_118_state = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  states_119_state = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  states_120_state = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  states_121_state = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  states_122_state = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  states_123_state = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  states_124_state = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  states_125_state = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  states_126_state = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  states_127_state = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  states_128_state = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  states_129_state = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  states_130_state = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  states_131_state = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  states_132_state = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  states_133_state = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  states_134_state = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  states_135_state = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  states_136_state = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  states_137_state = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  states_138_state = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  states_139_state = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  states_140_state = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  states_141_state = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  states_142_state = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  states_143_state = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  states_144_state = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  states_145_state = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  states_146_state = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  states_147_state = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  states_148_state = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  states_149_state = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  states_150_state = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  states_151_state = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  states_152_state = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  states_153_state = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  states_154_state = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  states_155_state = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  states_156_state = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  states_157_state = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  states_158_state = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  states_159_state = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  states_160_state = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  states_161_state = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  states_162_state = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  states_163_state = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  states_164_state = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  states_165_state = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  states_166_state = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  states_167_state = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  states_168_state = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  states_169_state = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  states_170_state = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  states_171_state = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  states_172_state = _RAND_172[1:0];
  _RAND_173 = {1{`RANDOM}};
  states_173_state = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  states_174_state = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  states_175_state = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  states_176_state = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  states_177_state = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  states_178_state = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  states_179_state = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  states_180_state = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  states_181_state = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  states_182_state = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  states_183_state = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  states_184_state = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  states_185_state = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  states_186_state = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  states_187_state = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  states_188_state = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  states_189_state = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  states_190_state = _RAND_190[1:0];
  _RAND_191 = {1{`RANDOM}};
  states_191_state = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  states_192_state = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  states_193_state = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  states_194_state = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  states_195_state = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  states_196_state = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  states_197_state = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  states_198_state = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  states_199_state = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  states_200_state = _RAND_200[1:0];
  _RAND_201 = {1{`RANDOM}};
  states_201_state = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  states_202_state = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  states_203_state = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  states_204_state = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  states_205_state = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  states_206_state = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  states_207_state = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  states_208_state = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  states_209_state = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  states_210_state = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  states_211_state = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  states_212_state = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  states_213_state = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  states_214_state = _RAND_214[1:0];
  _RAND_215 = {1{`RANDOM}};
  states_215_state = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  states_216_state = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  states_217_state = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  states_218_state = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  states_219_state = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  states_220_state = _RAND_220[1:0];
  _RAND_221 = {1{`RANDOM}};
  states_221_state = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  states_222_state = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  states_223_state = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  states_224_state = _RAND_224[1:0];
  _RAND_225 = {1{`RANDOM}};
  states_225_state = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  states_226_state = _RAND_226[1:0];
  _RAND_227 = {1{`RANDOM}};
  states_227_state = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  states_228_state = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  states_229_state = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  states_230_state = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  states_231_state = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  states_232_state = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  states_233_state = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  states_234_state = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  states_235_state = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  states_236_state = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  states_237_state = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  states_238_state = _RAND_238[1:0];
  _RAND_239 = {1{`RANDOM}};
  states_239_state = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  states_240_state = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  states_241_state = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  states_242_state = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  states_243_state = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  states_244_state = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  states_245_state = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  states_246_state = _RAND_246[1:0];
  _RAND_247 = {1{`RANDOM}};
  states_247_state = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  states_248_state = _RAND_248[1:0];
  _RAND_249 = {1{`RANDOM}};
  states_249_state = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  states_250_state = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  states_251_state = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  states_252_state = _RAND_252[1:0];
  _RAND_253 = {1{`RANDOM}};
  states_253_state = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  states_254_state = _RAND_254[1:0];
  _RAND_255 = {1{`RANDOM}};
  states_255_state = _RAND_255[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      states_0_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h0 == idxSet_0) begin
        states_0_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_1_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h1 == idxSet_0) begin
        states_1_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_2_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h2 == idxSet_0) begin
        states_2_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_3_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h3 == idxSet_0) begin
        states_3_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_4_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h4 == idxSet_0) begin
        states_4_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_5_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h5 == idxSet_0) begin
        states_5_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_6_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h6 == idxSet_0) begin
        states_6_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_7_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h7 == idxSet_0) begin
        states_7_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_8_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h8 == idxSet_0) begin
        states_8_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_9_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h9 == idxSet_0) begin
        states_9_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_10_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'ha == idxSet_0) begin
        states_10_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_11_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hb == idxSet_0) begin
        states_11_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_12_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hc == idxSet_0) begin
        states_12_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_13_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hd == idxSet_0) begin
        states_13_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_14_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'he == idxSet_0) begin
        states_14_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_15_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hf == idxSet_0) begin
        states_15_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_16_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h10 == idxSet_0) begin
        states_16_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_17_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h11 == idxSet_0) begin
        states_17_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_18_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h12 == idxSet_0) begin
        states_18_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_19_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h13 == idxSet_0) begin
        states_19_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_20_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h14 == idxSet_0) begin
        states_20_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_21_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h15 == idxSet_0) begin
        states_21_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_22_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h16 == idxSet_0) begin
        states_22_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_23_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h17 == idxSet_0) begin
        states_23_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_24_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h18 == idxSet_0) begin
        states_24_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_25_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h19 == idxSet_0) begin
        states_25_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_26_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h1a == idxSet_0) begin
        states_26_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_27_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h1b == idxSet_0) begin
        states_27_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_28_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h1c == idxSet_0) begin
        states_28_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_29_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h1d == idxSet_0) begin
        states_29_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_30_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h1e == idxSet_0) begin
        states_30_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_31_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h1f == idxSet_0) begin
        states_31_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_32_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h20 == idxSet_0) begin
        states_32_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_33_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h21 == idxSet_0) begin
        states_33_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_34_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h22 == idxSet_0) begin
        states_34_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_35_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h23 == idxSet_0) begin
        states_35_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_36_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h24 == idxSet_0) begin
        states_36_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_37_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h25 == idxSet_0) begin
        states_37_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_38_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h26 == idxSet_0) begin
        states_38_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_39_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h27 == idxSet_0) begin
        states_39_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_40_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h28 == idxSet_0) begin
        states_40_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_41_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h29 == idxSet_0) begin
        states_41_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_42_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h2a == idxSet_0) begin
        states_42_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_43_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h2b == idxSet_0) begin
        states_43_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_44_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h2c == idxSet_0) begin
        states_44_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_45_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h2d == idxSet_0) begin
        states_45_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_46_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h2e == idxSet_0) begin
        states_46_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_47_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h2f == idxSet_0) begin
        states_47_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_48_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h30 == idxSet_0) begin
        states_48_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_49_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h31 == idxSet_0) begin
        states_49_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_50_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h32 == idxSet_0) begin
        states_50_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_51_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h33 == idxSet_0) begin
        states_51_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_52_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h34 == idxSet_0) begin
        states_52_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_53_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h35 == idxSet_0) begin
        states_53_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_54_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h36 == idxSet_0) begin
        states_54_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_55_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h37 == idxSet_0) begin
        states_55_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_56_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h38 == idxSet_0) begin
        states_56_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_57_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h39 == idxSet_0) begin
        states_57_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_58_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h3a == idxSet_0) begin
        states_58_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_59_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h3b == idxSet_0) begin
        states_59_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_60_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h3c == idxSet_0) begin
        states_60_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_61_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h3d == idxSet_0) begin
        states_61_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_62_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h3e == idxSet_0) begin
        states_62_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_63_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h3f == idxSet_0) begin
        states_63_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_64_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h40 == idxSet_0) begin
        states_64_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_65_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h41 == idxSet_0) begin
        states_65_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_66_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h42 == idxSet_0) begin
        states_66_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_67_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h43 == idxSet_0) begin
        states_67_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_68_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h44 == idxSet_0) begin
        states_68_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_69_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h45 == idxSet_0) begin
        states_69_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_70_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h46 == idxSet_0) begin
        states_70_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_71_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h47 == idxSet_0) begin
        states_71_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_72_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h48 == idxSet_0) begin
        states_72_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_73_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h49 == idxSet_0) begin
        states_73_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_74_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h4a == idxSet_0) begin
        states_74_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_75_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h4b == idxSet_0) begin
        states_75_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_76_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h4c == idxSet_0) begin
        states_76_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_77_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h4d == idxSet_0) begin
        states_77_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_78_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h4e == idxSet_0) begin
        states_78_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_79_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h4f == idxSet_0) begin
        states_79_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_80_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h50 == idxSet_0) begin
        states_80_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_81_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h51 == idxSet_0) begin
        states_81_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_82_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h52 == idxSet_0) begin
        states_82_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_83_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h53 == idxSet_0) begin
        states_83_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_84_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h54 == idxSet_0) begin
        states_84_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_85_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h55 == idxSet_0) begin
        states_85_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_86_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h56 == idxSet_0) begin
        states_86_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_87_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h57 == idxSet_0) begin
        states_87_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_88_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h58 == idxSet_0) begin
        states_88_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_89_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h59 == idxSet_0) begin
        states_89_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_90_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h5a == idxSet_0) begin
        states_90_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_91_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h5b == idxSet_0) begin
        states_91_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_92_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h5c == idxSet_0) begin
        states_92_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_93_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h5d == idxSet_0) begin
        states_93_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_94_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h5e == idxSet_0) begin
        states_94_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_95_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h5f == idxSet_0) begin
        states_95_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_96_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h60 == idxSet_0) begin
        states_96_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_97_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h61 == idxSet_0) begin
        states_97_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_98_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h62 == idxSet_0) begin
        states_98_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_99_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h63 == idxSet_0) begin
        states_99_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_100_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h64 == idxSet_0) begin
        states_100_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_101_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h65 == idxSet_0) begin
        states_101_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_102_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h66 == idxSet_0) begin
        states_102_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_103_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h67 == idxSet_0) begin
        states_103_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_104_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h68 == idxSet_0) begin
        states_104_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_105_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h69 == idxSet_0) begin
        states_105_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_106_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h6a == idxSet_0) begin
        states_106_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_107_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h6b == idxSet_0) begin
        states_107_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_108_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h6c == idxSet_0) begin
        states_108_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_109_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h6d == idxSet_0) begin
        states_109_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_110_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h6e == idxSet_0) begin
        states_110_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_111_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h6f == idxSet_0) begin
        states_111_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_112_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h70 == idxSet_0) begin
        states_112_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_113_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h71 == idxSet_0) begin
        states_113_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_114_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h72 == idxSet_0) begin
        states_114_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_115_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h73 == idxSet_0) begin
        states_115_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_116_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h74 == idxSet_0) begin
        states_116_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_117_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h75 == idxSet_0) begin
        states_117_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_118_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h76 == idxSet_0) begin
        states_118_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_119_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h77 == idxSet_0) begin
        states_119_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_120_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h78 == idxSet_0) begin
        states_120_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_121_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h79 == idxSet_0) begin
        states_121_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_122_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h7a == idxSet_0) begin
        states_122_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_123_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h7b == idxSet_0) begin
        states_123_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_124_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h7c == idxSet_0) begin
        states_124_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_125_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h7d == idxSet_0) begin
        states_125_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_126_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h7e == idxSet_0) begin
        states_126_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_127_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h7f == idxSet_0) begin
        states_127_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_128_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h80 == idxSet_0) begin
        states_128_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_129_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h81 == idxSet_0) begin
        states_129_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_130_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h82 == idxSet_0) begin
        states_130_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_131_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h83 == idxSet_0) begin
        states_131_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_132_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h84 == idxSet_0) begin
        states_132_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_133_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h85 == idxSet_0) begin
        states_133_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_134_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h86 == idxSet_0) begin
        states_134_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_135_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h87 == idxSet_0) begin
        states_135_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_136_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h88 == idxSet_0) begin
        states_136_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_137_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h89 == idxSet_0) begin
        states_137_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_138_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h8a == idxSet_0) begin
        states_138_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_139_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h8b == idxSet_0) begin
        states_139_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_140_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h8c == idxSet_0) begin
        states_140_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_141_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h8d == idxSet_0) begin
        states_141_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_142_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h8e == idxSet_0) begin
        states_142_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_143_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h8f == idxSet_0) begin
        states_143_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_144_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h90 == idxSet_0) begin
        states_144_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_145_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h91 == idxSet_0) begin
        states_145_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_146_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h92 == idxSet_0) begin
        states_146_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_147_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h93 == idxSet_0) begin
        states_147_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_148_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h94 == idxSet_0) begin
        states_148_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_149_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h95 == idxSet_0) begin
        states_149_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_150_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h96 == idxSet_0) begin
        states_150_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_151_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h97 == idxSet_0) begin
        states_151_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_152_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h98 == idxSet_0) begin
        states_152_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_153_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h99 == idxSet_0) begin
        states_153_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_154_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h9a == idxSet_0) begin
        states_154_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_155_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h9b == idxSet_0) begin
        states_155_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_156_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h9c == idxSet_0) begin
        states_156_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_157_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h9d == idxSet_0) begin
        states_157_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_158_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h9e == idxSet_0) begin
        states_158_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_159_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'h9f == idxSet_0) begin
        states_159_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_160_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'ha0 == idxSet_0) begin
        states_160_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_161_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'ha1 == idxSet_0) begin
        states_161_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_162_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'ha2 == idxSet_0) begin
        states_162_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_163_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'ha3 == idxSet_0) begin
        states_163_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_164_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'ha4 == idxSet_0) begin
        states_164_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_165_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'ha5 == idxSet_0) begin
        states_165_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_166_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'ha6 == idxSet_0) begin
        states_166_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_167_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'ha7 == idxSet_0) begin
        states_167_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_168_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'ha8 == idxSet_0) begin
        states_168_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_169_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'ha9 == idxSet_0) begin
        states_169_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_170_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'haa == idxSet_0) begin
        states_170_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_171_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hab == idxSet_0) begin
        states_171_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_172_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hac == idxSet_0) begin
        states_172_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_173_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'had == idxSet_0) begin
        states_173_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_174_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hae == idxSet_0) begin
        states_174_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_175_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'haf == idxSet_0) begin
        states_175_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_176_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hb0 == idxSet_0) begin
        states_176_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_177_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hb1 == idxSet_0) begin
        states_177_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_178_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hb2 == idxSet_0) begin
        states_178_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_179_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hb3 == idxSet_0) begin
        states_179_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_180_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hb4 == idxSet_0) begin
        states_180_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_181_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hb5 == idxSet_0) begin
        states_181_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_182_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hb6 == idxSet_0) begin
        states_182_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_183_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hb7 == idxSet_0) begin
        states_183_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_184_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hb8 == idxSet_0) begin
        states_184_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_185_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hb9 == idxSet_0) begin
        states_185_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_186_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hba == idxSet_0) begin
        states_186_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_187_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hbb == idxSet_0) begin
        states_187_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_188_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hbc == idxSet_0) begin
        states_188_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_189_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hbd == idxSet_0) begin
        states_189_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_190_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hbe == idxSet_0) begin
        states_190_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_191_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hbf == idxSet_0) begin
        states_191_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_192_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hc0 == idxSet_0) begin
        states_192_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_193_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hc1 == idxSet_0) begin
        states_193_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_194_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hc2 == idxSet_0) begin
        states_194_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_195_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hc3 == idxSet_0) begin
        states_195_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_196_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hc4 == idxSet_0) begin
        states_196_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_197_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hc5 == idxSet_0) begin
        states_197_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_198_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hc6 == idxSet_0) begin
        states_198_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_199_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hc7 == idxSet_0) begin
        states_199_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_200_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hc8 == idxSet_0) begin
        states_200_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_201_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hc9 == idxSet_0) begin
        states_201_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_202_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hca == idxSet_0) begin
        states_202_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_203_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hcb == idxSet_0) begin
        states_203_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_204_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hcc == idxSet_0) begin
        states_204_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_205_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hcd == idxSet_0) begin
        states_205_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_206_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hce == idxSet_0) begin
        states_206_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_207_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hcf == idxSet_0) begin
        states_207_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_208_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hd0 == idxSet_0) begin
        states_208_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_209_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hd1 == idxSet_0) begin
        states_209_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_210_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hd2 == idxSet_0) begin
        states_210_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_211_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hd3 == idxSet_0) begin
        states_211_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_212_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hd4 == idxSet_0) begin
        states_212_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_213_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hd5 == idxSet_0) begin
        states_213_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_214_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hd6 == idxSet_0) begin
        states_214_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_215_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hd7 == idxSet_0) begin
        states_215_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_216_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hd8 == idxSet_0) begin
        states_216_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_217_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hd9 == idxSet_0) begin
        states_217_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_218_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hda == idxSet_0) begin
        states_218_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_219_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hdb == idxSet_0) begin
        states_219_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_220_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hdc == idxSet_0) begin
        states_220_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_221_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hdd == idxSet_0) begin
        states_221_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_222_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hde == idxSet_0) begin
        states_222_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_223_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hdf == idxSet_0) begin
        states_223_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_224_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'he0 == idxSet_0) begin
        states_224_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_225_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'he1 == idxSet_0) begin
        states_225_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_226_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'he2 == idxSet_0) begin
        states_226_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_227_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'he3 == idxSet_0) begin
        states_227_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_228_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'he4 == idxSet_0) begin
        states_228_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_229_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'he5 == idxSet_0) begin
        states_229_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_230_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'he6 == idxSet_0) begin
        states_230_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_231_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'he7 == idxSet_0) begin
        states_231_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_232_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'he8 == idxSet_0) begin
        states_232_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_233_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'he9 == idxSet_0) begin
        states_233_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_234_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hea == idxSet_0) begin
        states_234_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_235_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'heb == idxSet_0) begin
        states_235_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_236_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hec == idxSet_0) begin
        states_236_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_237_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hed == idxSet_0) begin
        states_237_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_238_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hee == idxSet_0) begin
        states_238_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_239_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hef == idxSet_0) begin
        states_239_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_240_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hf0 == idxSet_0) begin
        states_240_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_241_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hf1 == idxSet_0) begin
        states_241_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_242_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hf2 == idxSet_0) begin
        states_242_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_243_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hf3 == idxSet_0) begin
        states_243_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_244_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hf4 == idxSet_0) begin
        states_244_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_245_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hf5 == idxSet_0) begin
        states_245_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_246_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hf6 == idxSet_0) begin
        states_246_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_247_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hf7 == idxSet_0) begin
        states_247_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_248_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hf8 == idxSet_0) begin
        states_248_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_249_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hf9 == idxSet_0) begin
        states_249_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_250_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hfa == idxSet_0) begin
        states_250_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_251_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hfb == idxSet_0) begin
        states_251_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_252_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hfc == idxSet_0) begin
        states_252_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_253_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hfd == idxSet_0) begin
        states_253_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_254_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hfe == idxSet_0) begin
        states_254_state <= io_in_0_bits_state_state;
      end
    end
    if (reset) begin
      states_255_state <= 2'h0;
    end else if (isSet_0) begin
      if (8'hff == idxSet_0) begin
        states_255_state <= io_in_0_bits_state_state;
      end
    end
  end
endmodule
module FindEmptyLine_3(
  input   io_data_0,
  output  io_value_valid,
  output  io_value_bits
);
  wire  _T = ~io_data_0; // @[elements.scala 74:53]
  wire [1:0] idx = _T ? 2'h0 : 2'h1; // @[elements.scala 74:66]
  assign io_value_valid = ~io_data_0; // @[elements.scala 68:20 elements.scala 76:32]
  assign io_value_bits = idx[0]; // @[elements.scala 79:19]
endmodule
module PC(
  input         clock,
  input         reset,
  output        io_write_ready,
  input         io_write_valid,
  input  [31:0] io_write_bits_addr,
  input  [2:0]  io_write_bits_way,
  input  [63:0] io_write_bits_data,
  input  [2:0]  io_write_bits_replaceWay,
  input  [31:0] io_write_bits_tbeFields_0,
  input  [15:0] io_write_bits_pc,
  input  [2:0]  io_read_0_in_bits_data_way,
  input  [15:0] io_read_0_in_bits_data_pc,
  input         io_read_0_in_bits_data_valid,
  output [31:0] io_read_0_out_bits_addr,
  output [2:0]  io_read_0_out_bits_way,
  output [63:0] io_read_0_out_bits_data,
  output [2:0]  io_read_0_out_bits_replaceWay,
  output [31:0] io_read_0_out_bits_tbeFields_0,
  output [15:0] io_read_0_out_bits_pc,
  output        io_read_0_out_bits_valid,
  output        io_isFull
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  findNewLine_io_data_0; // @[elements.scala 278:29]
  wire  findNewLine_io_value_valid; // @[elements.scala 278:29]
  wire  findNewLine_io_value_bits; // @[elements.scala 278:29]
  reg [31:0] pcContent_0_addr; // @[elements.scala 274:29]
  reg [2:0] pcContent_0_way; // @[elements.scala 274:29]
  reg [63:0] pcContent_0_data; // @[elements.scala 274:29]
  reg [2:0] pcContent_0_replaceWay; // @[elements.scala 274:29]
  reg [31:0] pcContent_0_tbeFields_0; // @[elements.scala 274:29]
  reg [15:0] pcContent_0_pc; // @[elements.scala 274:29]
  reg  pcContent_0_valid; // @[elements.scala 274:29]
  wire  write = io_write_ready & io_write_valid; // @[Decoupled.scala 40:37]
  wire  _T_113 = ~write; // @[elements.scala 288:14]
  wire  writeIdx = findNewLine_io_value_bits;
  wire  _T_115 = write & writeIdx; // @[elements.scala 288:30]
  wire  _T_116 = _T_113 | _T_115; // @[elements.scala 288:21]
  wire  _GEN_1 = _T_116 ? io_read_0_in_bits_data_valid : pcContent_0_valid; // @[elements.scala 288:50]
  wire  _GEN_10 = write | _GEN_1; // @[elements.scala 295:17]
  FindEmptyLine_3 findNewLine ( // @[elements.scala 278:29]
    .io_data_0(findNewLine_io_data_0),
    .io_value_valid(findNewLine_io_value_valid),
    .io_value_bits(findNewLine_io_value_bits)
  );
  assign io_write_ready = findNewLine_io_value_valid; // @[elements.scala 299:20]
  assign io_read_0_out_bits_addr = pcContent_0_addr; // @[elements.scala 283:30]
  assign io_read_0_out_bits_way = pcContent_0_way; // @[elements.scala 283:30]
  assign io_read_0_out_bits_data = pcContent_0_data; // @[elements.scala 283:30]
  assign io_read_0_out_bits_replaceWay = pcContent_0_replaceWay; // @[elements.scala 283:30]
  assign io_read_0_out_bits_tbeFields_0 = pcContent_0_tbeFields_0; // @[elements.scala 283:30]
  assign io_read_0_out_bits_pc = pcContent_0_pc; // @[elements.scala 283:30]
  assign io_read_0_out_bits_valid = pcContent_0_valid; // @[elements.scala 283:30]
  assign io_isFull = ~io_write_ready; // @[elements.scala 300:15]
  assign findNewLine_io_data_0 = pcContent_0_valid; // @[elements.scala 279:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pcContent_0_addr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  pcContent_0_way = _RAND_1[2:0];
  _RAND_2 = {2{`RANDOM}};
  pcContent_0_data = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  pcContent_0_replaceWay = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  pcContent_0_tbeFields_0 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  pcContent_0_pc = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  pcContent_0_valid = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pcContent_0_addr <= 32'h0;
    end else if (write) begin
      pcContent_0_addr <= io_write_bits_addr;
    end
    if (reset) begin
      pcContent_0_way <= 3'h4;
    end else if (write) begin
      pcContent_0_way <= io_write_bits_way;
    end else if (_T_116) begin
      pcContent_0_way <= io_read_0_in_bits_data_way;
    end
    if (reset) begin
      pcContent_0_data <= 64'h0;
    end else if (write) begin
      pcContent_0_data <= io_write_bits_data;
    end
    if (reset) begin
      pcContent_0_replaceWay <= 3'h0;
    end else if (write) begin
      pcContent_0_replaceWay <= io_write_bits_replaceWay;
    end
    if (reset) begin
      pcContent_0_tbeFields_0 <= 32'h0;
    end else if (write) begin
      pcContent_0_tbeFields_0 <= io_write_bits_tbeFields_0;
    end
    if (reset) begin
      pcContent_0_pc <= 16'h0;
    end else if (write) begin
      pcContent_0_pc <= io_write_bits_pc;
    end else if (_T_116) begin
      pcContent_0_pc <= io_read_0_in_bits_data_pc;
    end
    if (reset) begin
      pcContent_0_valid <= 1'h0;
    end else begin
      pcContent_0_valid <= _GEN_10;
    end
  end
endmodule
module Arbiter_3(
  input         io_in_0_valid,
  input  [1:0]  io_in_0_bits_event,
  input  [31:0] io_in_0_bits_addr,
  input  [63:0] io_in_0_bits_data,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [1:0]  io_in_1_bits_event,
  input  [31:0] io_in_1_bits_addr,
  input  [63:0] io_in_1_bits_data,
  input         io_in_2_valid,
  input  [1:0]  io_in_2_bits_event,
  input  [31:0] io_in_2_bits_addr,
  input  [63:0] io_in_2_bits_data,
  input         io_in_3_valid,
  input  [1:0]  io_in_3_bits_event,
  input  [31:0] io_in_3_bits_addr,
  input  [63:0] io_in_3_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output [1:0]  io_out_bits_event,
  output [31:0] io_out_bits_addr,
  output [63:0] io_out_bits_data,
  output [1:0]  io_chosen
);
  wire [1:0] _GEN_0 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_1 = io_in_2_valid ? io_in_2_bits_data : io_in_3_bits_data; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_2 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_3 = io_in_2_valid ? io_in_2_bits_event : io_in_3_bits_event; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_4 = io_in_1_valid ? 2'h1 : _GEN_0; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_5 = io_in_1_valid ? io_in_1_bits_data : _GEN_1; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_6 = io_in_1_valid ? io_in_1_bits_addr : _GEN_2; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_7 = io_in_1_valid ? io_in_1_bits_event : _GEN_3; // @[Arbiter.scala 126:27]
  wire  _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  _T_1 = _T | io_in_2_valid; // @[Arbiter.scala 31:68]
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  grant_3 = ~_T_1; // @[Arbiter.scala 31:78]
  wire  _T_6 = ~grant_3; // @[Arbiter.scala 135:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_6 | io_in_3_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_event = io_in_0_valid ? io_in_0_bits_event : _GEN_7; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_6; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : _GEN_5; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_chosen = io_in_0_valid ? 2'h0 : _GEN_4; // @[Arbiter.scala 123:13 Arbiter.scala 127:17 Arbiter.scala 127:17 Arbiter.scala 127:17]
endmodule
module RRArbiter_2(
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_req_addr,
  input  [7:0]  io_in_0_bits_req_inst,
  input  [63:0] io_in_0_bits_req_data,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [7:0]  io_out_bits_req_inst,
  output [63:0] io_out_bits_req_data
);
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_req_addr = io_in_0_bits_req_addr; // @[Arbiter.scala 42:15]
  assign io_out_bits_req_inst = io_in_0_bits_req_inst; // @[Arbiter.scala 42:15]
  assign io_out_bits_req_data = io_in_0_bits_req_data; // @[Arbiter.scala 42:15]
endmodule
module Arbiter_4(
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  output        io_out_valid,
  output [31:0] io_out_bits_addr
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module Arbiter_5(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [1:0]  io_in_0_bits_event,
  input  [31:0] io_in_0_bits_addr,
  input  [63:0] io_in_0_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output [1:0]  io_out_bits_event,
  output [31:0] io_out_bits_addr,
  output [63:0] io_out_bits_data
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_event = io_in_0_bits_event; // @[Arbiter.scala 124:15]
  assign io_out_bits_addr = io_in_0_bits_addr; // @[Arbiter.scala 124:15]
  assign io_out_bits_data = io_in_0_bits_data; // @[Arbiter.scala 124:15]
endmodule
module Queue_7(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_inst_event,
  input  [31:0] io_enq_bits_inst_addr,
  input  [63:0] io_enq_bits_inst_data,
  input  [1:0]  io_enq_bits_tbeOut_state_state,
  input  [3:0]  io_enq_bits_tbeOut_way,
  input  [31:0] io_enq_bits_tbeOut_fields_0,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_inst_event,
  output [31:0] io_deq_bits_inst_addr,
  output [63:0] io_deq_bits_inst_data,
  output [1:0]  io_deq_bits_tbeOut_state_state,
  output [3:0]  io_deq_bits_tbeOut_way,
  output [31:0] io_deq_bits_tbeOut_fields_0
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_inst_event [0:0]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_inst_event__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_inst_event__T_7_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_inst_event__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst_event__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst_event__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst_event__T_3_en; // @[Decoupled.scala 209:16]
  reg [31:0] ram_inst_addr [0:0]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_inst_addr__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_inst_addr__T_7_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_inst_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_inst_data [0:0]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_inst_data__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_inst_data__T_7_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_inst_data__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [1:0] ram_tbeOut_state_state [0:0]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_tbeOut_state_state__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_state_state__T_7_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_tbeOut_state_state__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_state_state__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_state_state__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_state_state__T_3_en; // @[Decoupled.scala 209:16]
  reg [3:0] ram_tbeOut_way [0:0]; // @[Decoupled.scala 209:16]
  wire [3:0] ram_tbeOut_way__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_way__T_7_addr; // @[Decoupled.scala 209:16]
  wire [3:0] ram_tbeOut_way__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_way__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_way__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_way__T_3_en; // @[Decoupled.scala 209:16]
  reg [31:0] ram_tbeOut_fields_0 [0:0]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_tbeOut_fields_0__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_fields_0__T_7_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_tbeOut_fields_0__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_fields_0__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_fields_0__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_tbeOut_fields_0__T_3_en; // @[Decoupled.scala 209:16]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram_inst_event__T_7_addr = 1'h0;
  assign ram_inst_event__T_7_data = ram_inst_event[ram_inst_event__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst_event__T_3_data = io_enq_bits_inst_event;
  assign ram_inst_event__T_3_addr = 1'h0;
  assign ram_inst_event__T_3_mask = 1'h1;
  assign ram_inst_event__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst_addr__T_7_addr = 1'h0;
  assign ram_inst_addr__T_7_data = ram_inst_addr[ram_inst_addr__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst_addr__T_3_data = io_enq_bits_inst_addr;
  assign ram_inst_addr__T_3_addr = 1'h0;
  assign ram_inst_addr__T_3_mask = 1'h1;
  assign ram_inst_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst_data__T_7_addr = 1'h0;
  assign ram_inst_data__T_7_data = ram_inst_data[ram_inst_data__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst_data__T_3_data = io_enq_bits_inst_data;
  assign ram_inst_data__T_3_addr = 1'h0;
  assign ram_inst_data__T_3_mask = 1'h1;
  assign ram_inst_data__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_tbeOut_state_state__T_7_addr = 1'h0;
  assign ram_tbeOut_state_state__T_7_data = ram_tbeOut_state_state[ram_tbeOut_state_state__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_tbeOut_state_state__T_3_data = io_enq_bits_tbeOut_state_state;
  assign ram_tbeOut_state_state__T_3_addr = 1'h0;
  assign ram_tbeOut_state_state__T_3_mask = 1'h1;
  assign ram_tbeOut_state_state__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_tbeOut_way__T_7_addr = 1'h0;
  assign ram_tbeOut_way__T_7_data = ram_tbeOut_way[ram_tbeOut_way__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_tbeOut_way__T_3_data = io_enq_bits_tbeOut_way;
  assign ram_tbeOut_way__T_3_addr = 1'h0;
  assign ram_tbeOut_way__T_3_mask = 1'h1;
  assign ram_tbeOut_way__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_tbeOut_fields_0__T_7_addr = 1'h0;
  assign ram_tbeOut_fields_0__T_7_data = ram_tbeOut_fields_0[ram_tbeOut_fields_0__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_tbeOut_fields_0__T_3_data = io_enq_bits_tbeOut_fields_0;
  assign ram_tbeOut_fields_0__T_3_addr = 1'h0;
  assign ram_tbeOut_fields_0__T_3_mask = 1'h1;
  assign ram_tbeOut_fields_0__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_inst_event = ram_inst_event__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst_addr = ram_inst_addr__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst_data = ram_inst_data__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_tbeOut_state_state = ram_tbeOut_state_state__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_tbeOut_way = ram_tbeOut_way__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_tbeOut_fields_0 = ram_tbeOut_fields_0__T_7_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_inst_event[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_inst_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_inst_data[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tbeOut_state_state[initvar] = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tbeOut_way[initvar] = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tbeOut_fields_0[initvar] = _RAND_5[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  maybe_full = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_inst_event__T_3_en & ram_inst_event__T_3_mask) begin
      ram_inst_event[ram_inst_event__T_3_addr] <= ram_inst_event__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst_addr__T_3_en & ram_inst_addr__T_3_mask) begin
      ram_inst_addr[ram_inst_addr__T_3_addr] <= ram_inst_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst_data__T_3_en & ram_inst_data__T_3_mask) begin
      ram_inst_data[ram_inst_data__T_3_addr] <= ram_inst_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_tbeOut_state_state__T_3_en & ram_tbeOut_state_state__T_3_mask) begin
      ram_tbeOut_state_state[ram_tbeOut_state_state__T_3_addr] <= ram_tbeOut_state_state__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_tbeOut_way__T_3_en & ram_tbeOut_way__T_3_mask) begin
      ram_tbeOut_way[ram_tbeOut_way__T_3_addr] <= ram_tbeOut_way__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_tbeOut_fields_0__T_3_en & ram_tbeOut_fields_0__T_3_mask) begin
      ram_tbeOut_fields_0[ram_tbeOut_fields_0__T_3_addr] <= ram_tbeOut_fields_0__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_4) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_8(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_event,
  input  [31:0] io_enq_bits_addr,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_event,
  output [31:0] io_deq_bits_addr,
  output [63:0] io_deq_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_event [0:15]; // @[Decoupled.scala 209:16]
  wire [1:0] ram_event__T_11_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram_event__T_11_addr; // @[Decoupled.scala 209:16]
  wire [1:0] ram_event__T_3_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram_event__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_event__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_event__T_3_en; // @[Decoupled.scala 209:16]
  reg [31:0] ram_addr [0:15]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_11_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram_addr__T_11_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:15]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_11_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram_data__T_11_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 29:33]
  reg [3:0] deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _T_5 = enq_ptr_value + 4'h1; // @[Counter.scala 39:22]
  wire [3:0] _T_7 = deq_ptr_value + 4'h1; // @[Counter.scala 39:22]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  wire  _T_10 = ~full; // @[Decoupled.scala 232:19]
  assign ram_event__T_11_addr = deq_ptr_value;
  assign ram_event__T_11_data = ram_event[ram_event__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_event__T_3_data = io_enq_bits_event;
  assign ram_event__T_3_addr = enq_ptr_value;
  assign ram_event__T_3_mask = 1'h1;
  assign ram_event__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_addr__T_11_addr = deq_ptr_value;
  assign ram_addr__T_11_data = ram_addr[ram_addr__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_3_data = io_enq_bits_addr;
  assign ram_addr__T_3_addr = enq_ptr_value;
  assign ram_addr__T_3_mask = 1'h1;
  assign ram_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_11_addr = deq_ptr_value;
  assign ram_data__T_11_data = ram_data[ram_data__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = enq_ptr_value;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | _T_10; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_event = ram_event__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_addr = ram_addr__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_11_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_event[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_event__T_3_en & ram_event__T_3_mask) begin
      ram_event[ram_event__T_3_addr] <= ram_event__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_addr__T_3_en & ram_addr__T_3_mask) begin
      ram_addr[ram_addr__T_3_addr] <= ram_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 4'h0;
    end else if (do_enq) begin
      enq_ptr_value <= _T_5;
    end
    if (reset) begin
      deq_ptr_value <= 4'h0;
    end else if (do_deq) begin
      deq_ptr_value <= _T_7;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_10(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [63:0] io_enq_bits_data,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_inst,
  output [63:0] io_deq_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:31]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_11_data; // @[Decoupled.scala 209:16]
  wire [4:0] ram_addr__T_11_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire [4:0] ram_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [7:0] ram_inst [0:31]; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_11_data; // @[Decoupled.scala 209:16]
  wire [4:0] ram_inst__T_11_addr; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_3_data; // @[Decoupled.scala 209:16]
  wire [4:0] ram_inst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:31]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_11_data; // @[Decoupled.scala 209:16]
  wire [4:0] ram_data__T_11_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire [4:0] ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [4:0] enq_ptr_value; // @[Counter.scala 29:33]
  reg [4:0] deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire [4:0] _T_5 = enq_ptr_value + 5'h1; // @[Counter.scala 39:22]
  wire [4:0] _T_7 = deq_ptr_value + 5'h1; // @[Counter.scala 39:22]
  wire  _T_8 = do_enq != io_deq_valid; // @[Decoupled.scala 227:16]
  assign ram_addr__T_11_addr = deq_ptr_value;
  assign ram_addr__T_11_data = ram_addr[ram_addr__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_3_data = io_enq_bits_addr;
  assign ram_addr__T_3_addr = enq_ptr_value;
  assign ram_addr__T_3_mask = 1'h1;
  assign ram_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst__T_11_addr = deq_ptr_value;
  assign ram_inst__T_11_data = ram_inst[ram_inst__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst__T_3_data = 8'h0;
  assign ram_inst__T_3_addr = enq_ptr_value;
  assign ram_inst__T_3_mask = 1'h1;
  assign ram_inst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_11_addr = deq_ptr_value;
  assign ram_data__T_11_data = ram_data[ram_data__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = enq_ptr_value;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = 1'h1; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst = ram_inst__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_11_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram_inst[initvar] = _RAND_1[7:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_3_en & ram_addr__T_3_mask) begin
      ram_addr[ram_addr__T_3_addr] <= ram_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst__T_3_en & ram_inst__T_3_mask) begin
      ram_inst[ram_inst__T_3_addr] <= ram_inst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 5'h0;
    end else if (do_enq) begin
      enq_ptr_value <= _T_5;
    end
    if (reset) begin
      deq_ptr_value <= 5'h0;
    end else if (io_deq_valid) begin
      deq_ptr_value <= _T_7;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_12(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram [0:15]; // @[Decoupled.scala 209:16]
  wire [2:0] ram__T_11_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram__T_11_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram__T_3_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram__T_3_en; // @[Decoupled.scala 209:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 29:33]
  reg [3:0] deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  _T_1 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _T_5 = enq_ptr_value + 4'h1; // @[Counter.scala 39:22]
  wire  _GEN_9 = io_deq_ready ? 1'h0 : _T_1; // @[Decoupled.scala 240:27]
  wire  do_enq = empty ? _GEN_9 : _T_1; // @[Decoupled.scala 237:18]
  wire [3:0] _T_7 = deq_ptr_value + 4'h1; // @[Counter.scala 39:22]
  wire  do_deq = empty ? 1'h0 : _T_2; // @[Decoupled.scala 237:18]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  wire  _T_9 = ~empty; // @[Decoupled.scala 231:19]
  wire  _T_10 = ~full; // @[Decoupled.scala 232:19]
  assign ram__T_11_addr = deq_ptr_value;
  assign ram__T_11_data = ram[ram__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram__T_3_data = io_enq_bits;
  assign ram__T_3_addr = enq_ptr_value;
  assign ram__T_3_mask = 1'h1;
  assign ram__T_3_en = empty ? _GEN_9 : _T_1;
  assign io_enq_ready = io_deq_ready | _T_10; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = io_enq_valid | _T_9; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits = empty ? io_enq_bits : ram__T_11_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram[initvar] = _RAND_0[2:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_3_en & ram__T_3_mask) begin
      ram[ram__T_3_addr] <= ram__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 4'h0;
    end else if (do_enq) begin
      enq_ptr_value <= _T_5;
    end
    if (reset) begin
      deq_ptr_value <= 4'h0;
    end else if (do_deq) begin
      deq_ptr_value <= _T_7;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _T_1;
        end
      end else begin
        maybe_full <= _T_1;
      end
    end
  end
endmodule
module Queue_14(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] ram [0:0]; // @[Decoupled.scala 209:16]
  wire [15:0] ram__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram__T_7_addr; // @[Decoupled.scala 209:16]
  wire [15:0] ram__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram__T_3_en; // @[Decoupled.scala 209:16]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram__T_7_addr = 1'h0;
  assign ram__T_7_data = ram[ram__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram__T_3_data = io_enq_bits;
  assign ram__T_3_addr = 1'h0;
  assign ram__T_3_mask = 1'h1;
  assign ram__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits = ram__T_7_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maybe_full = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_3_en & ram__T_3_mask) begin
      ram[ram__T_3_addr] <= ram__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_4) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_15(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [2:0]  io_enq_bits_way,
  input  [63:0] io_enq_bits_data,
  input  [2:0]  io_enq_bits_replaceWay,
  input  [31:0] io_enq_bits_tbeFields_0,
  input  [27:0] io_enq_bits_action_signals,
  input  [3:0]  io_enq_bits_action_actionType,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [2:0]  io_deq_bits_way,
  output [63:0] io_deq_bits_data,
  output [2:0]  io_deq_bits_replaceWay,
  output [31:0] io_deq_bits_tbeFields_0,
  output [27:0] io_deq_bits_action_signals,
  output [3:0]  io_deq_bits_action_actionType
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:0]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_33_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_27_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_way [0:0]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_way__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_way__T_33_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_way__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_way__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_way__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_way__T_27_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:0]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_33_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_27_en; // @[Decoupled.scala 209:16]
  reg [2:0] ram_replaceWay [0:0]; // @[Decoupled.scala 209:16]
  wire [2:0] ram_replaceWay__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_replaceWay__T_33_addr; // @[Decoupled.scala 209:16]
  wire [2:0] ram_replaceWay__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_replaceWay__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_replaceWay__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_replaceWay__T_27_en; // @[Decoupled.scala 209:16]
  reg [31:0] ram_tbeFields_0 [0:0]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_tbeFields_0__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeFields_0__T_33_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_tbeFields_0__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_tbeFields_0__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_tbeFields_0__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_tbeFields_0__T_27_en; // @[Decoupled.scala 209:16]
  reg [27:0] ram_action_signals [0:0]; // @[Decoupled.scala 209:16]
  wire [27:0] ram_action_signals__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_action_signals__T_33_addr; // @[Decoupled.scala 209:16]
  wire [27:0] ram_action_signals__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_action_signals__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_action_signals__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_action_signals__T_27_en; // @[Decoupled.scala 209:16]
  reg [3:0] ram_action_actionType [0:0]; // @[Decoupled.scala 209:16]
  wire [3:0] ram_action_actionType__T_33_data; // @[Decoupled.scala 209:16]
  wire  ram_action_actionType__T_33_addr; // @[Decoupled.scala 209:16]
  wire [3:0] ram_action_actionType__T_27_data; // @[Decoupled.scala 209:16]
  wire  ram_action_actionType__T_27_addr; // @[Decoupled.scala 209:16]
  wire  ram_action_actionType__T_27_mask; // @[Decoupled.scala 209:16]
  wire  ram_action_actionType__T_27_en; // @[Decoupled.scala 209:16]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = do_enq != io_deq_valid; // @[Decoupled.scala 227:16]
  assign ram_addr__T_33_addr = 1'h0;
  assign ram_addr__T_33_data = ram_addr[ram_addr__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_27_data = io_enq_bits_addr;
  assign ram_addr__T_27_addr = 1'h0;
  assign ram_addr__T_27_mask = 1'h1;
  assign ram_addr__T_27_en = io_enq_ready & io_enq_valid;
  assign ram_way__T_33_addr = 1'h0;
  assign ram_way__T_33_data = ram_way[ram_way__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_way__T_27_data = io_enq_bits_way;
  assign ram_way__T_27_addr = 1'h0;
  assign ram_way__T_27_mask = 1'h1;
  assign ram_way__T_27_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_33_addr = 1'h0;
  assign ram_data__T_33_data = ram_data[ram_data__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_27_data = io_enq_bits_data;
  assign ram_data__T_27_addr = 1'h0;
  assign ram_data__T_27_mask = 1'h1;
  assign ram_data__T_27_en = io_enq_ready & io_enq_valid;
  assign ram_replaceWay__T_33_addr = 1'h0;
  assign ram_replaceWay__T_33_data = ram_replaceWay[ram_replaceWay__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_replaceWay__T_27_data = io_enq_bits_replaceWay;
  assign ram_replaceWay__T_27_addr = 1'h0;
  assign ram_replaceWay__T_27_mask = 1'h1;
  assign ram_replaceWay__T_27_en = io_enq_ready & io_enq_valid;
  assign ram_tbeFields_0__T_33_addr = 1'h0;
  assign ram_tbeFields_0__T_33_data = ram_tbeFields_0[ram_tbeFields_0__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_tbeFields_0__T_27_data = io_enq_bits_tbeFields_0;
  assign ram_tbeFields_0__T_27_addr = 1'h0;
  assign ram_tbeFields_0__T_27_mask = 1'h1;
  assign ram_tbeFields_0__T_27_en = io_enq_ready & io_enq_valid;
  assign ram_action_signals__T_33_addr = 1'h0;
  assign ram_action_signals__T_33_data = ram_action_signals[ram_action_signals__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_action_signals__T_27_data = io_enq_bits_action_signals;
  assign ram_action_signals__T_27_addr = 1'h0;
  assign ram_action_signals__T_27_mask = 1'h1;
  assign ram_action_signals__T_27_en = io_enq_ready & io_enq_valid;
  assign ram_action_actionType__T_33_addr = 1'h0;
  assign ram_action_actionType__T_33_data = ram_action_actionType[ram_action_actionType__T_33_addr]; // @[Decoupled.scala 209:16]
  assign ram_action_actionType__T_27_data = io_enq_bits_action_actionType;
  assign ram_action_actionType__T_27_addr = 1'h0;
  assign ram_action_actionType__T_27_mask = 1'h1;
  assign ram_action_actionType__T_27_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = 1'h1; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_33_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_way = ram_way__T_33_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_33_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_replaceWay = ram_replaceWay__T_33_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_tbeFields_0 = ram_tbeFields_0__T_33_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_action_signals = ram_action_signals__T_33_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_action_actionType = ram_action_actionType__T_33_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_way[initvar] = _RAND_1[2:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_replaceWay[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tbeFields_0[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_action_signals[initvar] = _RAND_5[27:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_action_actionType[initvar] = _RAND_6[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_27_en & ram_addr__T_27_mask) begin
      ram_addr[ram_addr__T_27_addr] <= ram_addr__T_27_data; // @[Decoupled.scala 209:16]
    end
    if(ram_way__T_27_en & ram_way__T_27_mask) begin
      ram_way[ram_way__T_27_addr] <= ram_way__T_27_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_27_en & ram_data__T_27_mask) begin
      ram_data[ram_data__T_27_addr] <= ram_data__T_27_data; // @[Decoupled.scala 209:16]
    end
    if(ram_replaceWay__T_27_en & ram_replaceWay__T_27_mask) begin
      ram_replaceWay[ram_replaceWay__T_27_addr] <= ram_replaceWay__T_27_data; // @[Decoupled.scala 209:16]
    end
    if(ram_tbeFields_0__T_27_en & ram_tbeFields_0__T_27_mask) begin
      ram_tbeFields_0[ram_tbeFields_0__T_27_addr] <= ram_tbeFields_0__T_27_data; // @[Decoupled.scala 209:16]
    end
    if(ram_action_signals__T_27_en & ram_action_signals__T_27_mask) begin
      ram_action_signals[ram_action_signals__T_27_addr] <= ram_action_signals__T_27_data; // @[Decoupled.scala 209:16]
    end
    if(ram_action_actionType__T_27_en & ram_action_actionType__T_27_mask) begin
      ram_action_actionType[ram_action_actionType__T_27_addr] <= ram_action_actionType__T_27_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_30) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module MIMOQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_0_way,
  input  [31:0] io_enq_bits_0_addr,
  input  [2:0]  io_enq_bits_1_way,
  input  [31:0] io_enq_bits_1_addr,
  input  [2:0]  io_enq_bits_2_way,
  input  [31:0] io_enq_bits_2_addr,
  input  [2:0]  io_enq_bits_3_way,
  input  [31:0] io_enq_bits_3_addr,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_0_way,
  output [31:0] io_deq_bits_0_addr,
  output [7:0]  io_count
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_way [0:127]; // @[MIMOQueue.scala 56:16]
  wire [2:0] ram_way__T_28_data; // @[MIMOQueue.scala 56:16]
  wire [6:0] ram_way__T_28_addr; // @[MIMOQueue.scala 56:16]
  wire [2:0] ram_way__T_7_data; // @[MIMOQueue.scala 56:16]
  wire [6:0] ram_way__T_7_addr; // @[MIMOQueue.scala 56:16]
  wire  ram_way__T_7_mask; // @[MIMOQueue.scala 56:16]
  wire  ram_way__T_7_en; // @[MIMOQueue.scala 56:16]
  wire [2:0] ram_way__T_10_data; // @[MIMOQueue.scala 56:16]
  wire [6:0] ram_way__T_10_addr; // @[MIMOQueue.scala 56:16]
  wire  ram_way__T_10_mask; // @[MIMOQueue.scala 56:16]
  wire  ram_way__T_10_en; // @[MIMOQueue.scala 56:16]
  wire [2:0] ram_way__T_13_data; // @[MIMOQueue.scala 56:16]
  wire [6:0] ram_way__T_13_addr; // @[MIMOQueue.scala 56:16]
  wire  ram_way__T_13_mask; // @[MIMOQueue.scala 56:16]
  wire  ram_way__T_13_en; // @[MIMOQueue.scala 56:16]
  wire [2:0] ram_way__T_16_data; // @[MIMOQueue.scala 56:16]
  wire [6:0] ram_way__T_16_addr; // @[MIMOQueue.scala 56:16]
  wire  ram_way__T_16_mask; // @[MIMOQueue.scala 56:16]
  wire  ram_way__T_16_en; // @[MIMOQueue.scala 56:16]
  reg [31:0] ram_addr [0:127]; // @[MIMOQueue.scala 56:16]
  wire [31:0] ram_addr__T_28_data; // @[MIMOQueue.scala 56:16]
  wire [6:0] ram_addr__T_28_addr; // @[MIMOQueue.scala 56:16]
  wire [31:0] ram_addr__T_7_data; // @[MIMOQueue.scala 56:16]
  wire [6:0] ram_addr__T_7_addr; // @[MIMOQueue.scala 56:16]
  wire  ram_addr__T_7_mask; // @[MIMOQueue.scala 56:16]
  wire  ram_addr__T_7_en; // @[MIMOQueue.scala 56:16]
  wire [31:0] ram_addr__T_10_data; // @[MIMOQueue.scala 56:16]
  wire [6:0] ram_addr__T_10_addr; // @[MIMOQueue.scala 56:16]
  wire  ram_addr__T_10_mask; // @[MIMOQueue.scala 56:16]
  wire  ram_addr__T_10_en; // @[MIMOQueue.scala 56:16]
  wire [31:0] ram_addr__T_13_data; // @[MIMOQueue.scala 56:16]
  wire [6:0] ram_addr__T_13_addr; // @[MIMOQueue.scala 56:16]
  wire  ram_addr__T_13_mask; // @[MIMOQueue.scala 56:16]
  wire  ram_addr__T_13_en; // @[MIMOQueue.scala 56:16]
  wire [31:0] ram_addr__T_16_data; // @[MIMOQueue.scala 56:16]
  wire [6:0] ram_addr__T_16_addr; // @[MIMOQueue.scala 56:16]
  wire  ram_addr__T_16_mask; // @[MIMOQueue.scala 56:16]
  wire  ram_addr__T_16_en; // @[MIMOQueue.scala 56:16]
  reg [6:0] value; // @[Counter.scala 29:33]
  reg [6:0] value_1; // @[Counter.scala 29:33]
  reg  maybe_full; // @[MIMOQueue.scala 59:27]
  wire  ptr_match = value == value_1; // @[MIMOQueue.scala 62:33]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire [7:0] _T_5 = {{1'd0}, value}; // @[MIMOQueue.scala 77:25]
  wire [6:0] _T_18 = value + 7'h4; // @[MIMOQueue.scala 79:36]
  wire [6:0] _T_20 = value_1 + 7'h1; // @[MIMOQueue.scala 86:36]
  wire  _T_21 = do_enq != io_deq_valid; // @[MIMOQueue.scala 91:16]
  wire [6:0] ptr_diff = value - value_1; // @[MIMOQueue.scala 97:32]
  wire  _T_24 = io_count > 8'h0; // @[MIMOQueue.scala 100:18]
  wire [7:0] _T_26 = {{1'd0}, value_1}; // @[MIMOQueue.scala 106:73]
  wire  _T_31 = maybe_full & ptr_match; // @[MIMOQueue.scala 123:32]
  assign ram_way__T_28_addr = _T_26[6:0];
  assign ram_way__T_28_data = ram_way[ram_way__T_28_addr]; // @[MIMOQueue.scala 56:16]
  assign ram_way__T_7_data = io_enq_bits_0_way;
  assign ram_way__T_7_addr = _T_5[6:0];
  assign ram_way__T_7_mask = 1'h1;
  assign ram_way__T_7_en = io_enq_ready & io_enq_valid;
  assign ram_way__T_10_data = io_enq_bits_1_way;
  assign ram_way__T_10_addr = value + 7'h1;
  assign ram_way__T_10_mask = 1'h1;
  assign ram_way__T_10_en = io_enq_ready & io_enq_valid;
  assign ram_way__T_13_data = io_enq_bits_2_way;
  assign ram_way__T_13_addr = value + 7'h2;
  assign ram_way__T_13_mask = 1'h1;
  assign ram_way__T_13_en = io_enq_ready & io_enq_valid;
  assign ram_way__T_16_data = io_enq_bits_3_way;
  assign ram_way__T_16_addr = value + 7'h3;
  assign ram_way__T_16_mask = 1'h1;
  assign ram_way__T_16_en = io_enq_ready & io_enq_valid;
  assign ram_addr__T_28_addr = _T_26[6:0];
  assign ram_addr__T_28_data = ram_addr[ram_addr__T_28_addr]; // @[MIMOQueue.scala 56:16]
  assign ram_addr__T_7_data = io_enq_bits_0_addr;
  assign ram_addr__T_7_addr = _T_5[6:0];
  assign ram_addr__T_7_mask = 1'h1;
  assign ram_addr__T_7_en = io_enq_ready & io_enq_valid;
  assign ram_addr__T_10_data = io_enq_bits_1_addr;
  assign ram_addr__T_10_addr = value + 7'h1;
  assign ram_addr__T_10_mask = 1'h1;
  assign ram_addr__T_10_en = io_enq_ready & io_enq_valid;
  assign ram_addr__T_13_data = io_enq_bits_2_addr;
  assign ram_addr__T_13_addr = value + 7'h2;
  assign ram_addr__T_13_mask = 1'h1;
  assign ram_addr__T_13_en = io_enq_ready & io_enq_valid;
  assign ram_addr__T_16_data = io_enq_bits_3_addr;
  assign ram_addr__T_16_addr = value + 7'h3;
  assign ram_addr__T_16_mask = 1'h1;
  assign ram_addr__T_16_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = 1'h1; // @[MIMOQueue.scala 95:16 MIMOQueue.scala 119:40]
  assign io_deq_valid = io_count > 8'h0; // @[MIMOQueue.scala 101:18 MIMOQueue.scala 103:18]
  assign io_deq_bits_0_way = _T_24 ? ram_way__T_28_data : 3'h0; // @[MIMOQueue.scala 106:20]
  assign io_deq_bits_0_addr = _T_24 ? ram_addr__T_28_data : 32'h0; // @[MIMOQueue.scala 106:20]
  assign io_count = _T_31 ? 8'h80 : {{1'd0}, ptr_diff}; // @[MIMOQueue.scala 123:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_way[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_way__T_7_en & ram_way__T_7_mask) begin
      ram_way[ram_way__T_7_addr] <= ram_way__T_7_data; // @[MIMOQueue.scala 56:16]
    end
    if(ram_way__T_10_en & ram_way__T_10_mask) begin
      ram_way[ram_way__T_10_addr] <= ram_way__T_10_data; // @[MIMOQueue.scala 56:16]
    end
    if(ram_way__T_13_en & ram_way__T_13_mask) begin
      ram_way[ram_way__T_13_addr] <= ram_way__T_13_data; // @[MIMOQueue.scala 56:16]
    end
    if(ram_way__T_16_en & ram_way__T_16_mask) begin
      ram_way[ram_way__T_16_addr] <= ram_way__T_16_data; // @[MIMOQueue.scala 56:16]
    end
    if(ram_addr__T_7_en & ram_addr__T_7_mask) begin
      ram_addr[ram_addr__T_7_addr] <= ram_addr__T_7_data; // @[MIMOQueue.scala 56:16]
    end
    if(ram_addr__T_10_en & ram_addr__T_10_mask) begin
      ram_addr[ram_addr__T_10_addr] <= ram_addr__T_10_data; // @[MIMOQueue.scala 56:16]
    end
    if(ram_addr__T_13_en & ram_addr__T_13_mask) begin
      ram_addr[ram_addr__T_13_addr] <= ram_addr__T_13_data; // @[MIMOQueue.scala 56:16]
    end
    if(ram_addr__T_16_en & ram_addr__T_16_mask) begin
      ram_addr[ram_addr__T_16_addr] <= ram_addr__T_16_data; // @[MIMOQueue.scala 56:16]
    end
    if (reset) begin
      value <= 7'h0;
    end else if (do_enq) begin
      value <= _T_18;
    end
    if (reset) begin
      value_1 <= 7'h0;
    end else if (io_deq_valid) begin
      value_1 <= _T_20;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_21) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Computation(
  input         clock,
  input         reset,
  input         io_instruction_valid,
  input  [27:0] io_instruction_bits,
  input         io_clear,
  input         io_op1_valid,
  input  [63:0] io_op1_bits,
  input         io_op2_valid,
  input  [63:0] io_op2_bits,
  output [15:0] io_pc,
  output [63:0] io_reg_file_0,
  output [63:0] io_reg_file_1,
  output [63:0] io_reg_file_2,
  output [63:0] io_reg_file_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] function_ = io_instruction_bits[3:0]; // @[Computation.scala 69:42]
  wire [5:0] write_addr = io_instruction_bits[9:4]; // @[Computation.scala 70:42]
  wire [1:0] read_addr1 = io_instruction_bits[11:10]; // @[Computation.scala 73:42]
  wire [15:0] read_addr2 = io_instruction_bits[27:12]; // @[Computation.scala 74:42]
  reg [63:0] reg_file_3; // @[Computation.scala 86:27]
  reg [63:0] reg_file_2; // @[Computation.scala 86:27]
  reg [63:0] reg_file_1; // @[Computation.scala 86:27]
  reg [63:0] reg_file_0; // @[Computation.scala 86:27]
  wire [63:0] _GEN_13 = 2'h1 == read_addr1 ? reg_file_1 : reg_file_0; // @[Computation.scala 92:14]
  wire [63:0] _GEN_14 = 2'h2 == read_addr1 ? reg_file_2 : _GEN_13; // @[Computation.scala 92:14]
  wire [63:0] reg_out1 = 2'h3 == read_addr1 ? reg_file_3 : _GEN_14; // @[Computation.scala 92:14]
  wire [63:0] alu_in1 = io_op1_valid ? io_op1_bits : reg_out1; // @[Computation.scala 82:19]
  wire [63:0] _GEN_17 = 2'h1 == read_addr2[1:0] ? reg_file_1 : reg_file_0; // @[Computation.scala 93:14]
  wire [63:0] _GEN_18 = 2'h2 == read_addr2[1:0] ? reg_file_2 : _GEN_17; // @[Computation.scala 93:14]
  wire [63:0] reg_out2 = 2'h3 == read_addr2[1:0] ? reg_file_3 : _GEN_18; // @[Computation.scala 93:14]
  wire [63:0] alu_in2 = io_op2_valid ? io_op2_bits : reg_out2; // @[Computation.scala 83:19]
  wire  _T_3 = function_ != 4'h6; // @[Computation.scala 88:55]
  wire  _T_4 = function_ != 4'h7; // @[Computation.scala 88:75]
  wire  _T_5 = _T_3 & _T_4; // @[Computation.scala 88:63]
  wire  write_en = io_instruction_valid & _T_5; // @[Computation.scala 88:42]
  wire  _T_10 = 4'h0 == function_; // @[Conditional.scala 37:30]
  wire [63:0] _T_12 = alu_in1 + alu_in2; // @[Computation.scala 33:38]
  wire  _T_13 = 4'h1 == function_; // @[Conditional.scala 37:30]
  wire [63:0] _T_14 = alu_in1 & alu_in2; // @[Computation.scala 34:38]
  wire  _T_15 = 4'h2 == function_; // @[Conditional.scala 37:30]
  wire [63:0] _T_17 = alu_in1 - alu_in2; // @[Computation.scala 35:38]
  wire  _T_18 = 4'h3 == function_; // @[Conditional.scala 37:30]
  wire [63:0] _T_19 = alu_in1 >> alu_in2; // @[Computation.scala 36:42]
  wire  _T_20 = 4'h4 == function_; // @[Conditional.scala 37:30]
  wire [318:0] _GEN_29 = {{255'd0}, alu_in1}; // @[Computation.scala 37:42]
  wire [318:0] _T_22 = _GEN_29 << alu_in2[7:0]; // @[Computation.scala 37:42]
  wire  _T_23 = 4'h5 == function_; // @[Conditional.scala 37:30]
  wire [63:0] _T_24 = alu_in1 ^ alu_in2; // @[Computation.scala 38:38]
  wire  _T_25 = 4'h6 == function_; // @[Conditional.scala 37:30]
  wire  _T_26 = alu_in1 < alu_in2; // @[Computation.scala 39:43]
  wire [63:0] _T_8 = {{58'd0}, write_addr}; // @[Computation.scala 97:93 Computation.scala 97:93]
  wire [63:0] _T_27 = _T_26 ? _T_8 : 64'h0; // @[Computation.scala 39:38]
  wire  _T_28 = 4'h7 == function_; // @[Conditional.scala 37:30]
  wire  _T_29 = alu_in1 != alu_in2; // @[Computation.scala 40:43]
  wire [63:0] _T_30 = _T_29 ? _T_8 : 64'h0; // @[Computation.scala 40:38]
  wire  _T_31 = 4'h8 == function_; // @[Conditional.scala 37:30]
  wire [63:0] _T_32 = alu_in1 | alu_in2; // @[Computation.scala 41:37]
  wire [63:0] _GEN_20 = _T_31 ? _T_32 : 64'h0; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_21 = _T_28 ? _T_30 : _GEN_20; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_22 = _T_25 ? _T_27 : _GEN_21; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_23 = _T_23 ? _T_24 : _GEN_22; // @[Conditional.scala 39:67]
  wire [318:0] _GEN_24 = _T_20 ? _T_22 : {{255'd0}, _GEN_23}; // @[Conditional.scala 39:67]
  wire [318:0] _GEN_25 = _T_18 ? {{255'd0}, _T_19} : _GEN_24; // @[Conditional.scala 39:67]
  wire [318:0] _GEN_26 = _T_15 ? {{255'd0}, _T_17} : _GEN_25; // @[Conditional.scala 39:67]
  wire [318:0] _GEN_27 = _T_13 ? {{255'd0}, _T_14} : _GEN_26; // @[Conditional.scala 39:67]
  wire [318:0] _GEN_28 = _T_10 ? {{255'd0}, _T_12} : _GEN_27; // @[Conditional.scala 40:58]
  wire [63:0] result = io_instruction_valid ? _GEN_28[63:0] : 64'h0; // @[Computation.scala 97:18]
  assign io_pc = _T_5 ? 16'h0 : result[15:0]; // @[Computation.scala 98:11]
  assign io_reg_file_0 = reg_file_0; // @[Computation.scala 94:17]
  assign io_reg_file_1 = reg_file_1; // @[Computation.scala 94:17]
  assign io_reg_file_2 = reg_file_2; // @[Computation.scala 94:17]
  assign io_reg_file_3 = reg_file_3; // @[Computation.scala 94:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  reg_file_3 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  reg_file_2 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  reg_file_1 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  reg_file_0 = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      reg_file_3 <= 64'h0;
    end else if (io_clear) begin
      reg_file_3 <= 64'h0;
    end else if (write_en) begin
      if (2'h3 == write_addr[1:0]) begin
        if (io_instruction_valid) begin
          reg_file_3 <= _GEN_28[63:0];
        end else begin
          reg_file_3 <= 64'h0;
        end
      end
    end
    if (reset) begin
      reg_file_2 <= 64'h0;
    end else if (io_clear) begin
      reg_file_2 <= 64'h0;
    end else if (write_en) begin
      if (2'h2 == write_addr[1:0]) begin
        if (io_instruction_valid) begin
          reg_file_2 <= _GEN_28[63:0];
        end else begin
          reg_file_2 <= 64'h0;
        end
      end
    end
    if (reset) begin
      reg_file_1 <= 64'h0;
    end else if (io_clear) begin
      reg_file_1 <= 64'h0;
    end else if (write_en) begin
      if (2'h1 == write_addr[1:0]) begin
        if (io_instruction_valid) begin
          reg_file_1 <= _GEN_28[63:0];
        end else begin
          reg_file_1 <= 64'h0;
        end
      end
    end
    if (reset) begin
      reg_file_0 <= 64'h0;
    end else if (io_clear) begin
      reg_file_0 <= 64'h0;
    end else if (write_en) begin
      if (2'h0 == write_addr[1:0]) begin
        if (io_instruction_valid) begin
          reg_file_0 <= _GEN_28[63:0];
        end else begin
          reg_file_0 <= 64'h0;
        end
      end
    end
  end
endmodule
module Mux3(
  input  [63:0] io_in_hardCoded,
  input  [63:0] io_in_data,
  input  [63:0] io_in_tbe,
  input  [1:0]  io_in_select,
  output        io_out_valid,
  output [63:0] io_out_bits
);
  wire  _T = io_in_select == 2'h3; // @[ComputationUtils.scala 27:24]
  wire  _T_1 = io_in_select == 2'h2; // @[ComputationUtils.scala 29:31]
  wire  _T_2 = io_in_select == 2'h1; // @[ComputationUtils.scala 31:31]
  wire [63:0] _GEN_0 = _T_2 ? io_in_tbe : 64'h0; // @[ComputationUtils.scala 31:40]
  wire [63:0] _GEN_1 = _T_1 ? io_in_data : _GEN_0; // @[ComputationUtils.scala 29:40]
  wire [63:0] result = _T ? io_in_hardCoded : _GEN_1; // @[ComputationUtils.scala 27:33]
  assign io_out_valid = result != 64'h0; // @[ComputationUtils.scala 38:18]
  assign io_out_bits = _T ? io_in_hardCoded : _GEN_1; // @[ComputationUtils.scala 37:17]
endmodule
module programmableCache(
  input         clock,
  input         reset,
  output        io_in_cpu_ready,
  input         io_in_cpu_valid,
  input  [1:0]  io_in_cpu_bits_event,
  input  [31:0] io_in_cpu_bits_addr,
  input  [63:0] io_in_cpu_bits_data,
  output        io_in_memCtrl_ready,
  input         io_in_memCtrl_valid,
  input  [1:0]  io_in_memCtrl_bits_event,
  input  [31:0] io_in_memCtrl_bits_addr,
  input  [63:0] io_in_memCtrl_bits_data,
  output        io_in_otherNodes_ready,
  input         io_in_otherNodes_valid,
  input  [1:0]  io_in_otherNodes_bits_event,
  input  [31:0] io_in_otherNodes_bits_addr,
  input  [63:0] io_in_otherNodes_bits_data,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_req_addr,
  output [7:0]  io_out_req_bits_req_inst,
  output [63:0] io_out_req_bits_req_data,
  output        io_out_resp_valid,
  output [31:0] io_out_resp_bits_addr,
  output        _T_297_0,
  output        _T_291_0,
  output        _T_304_0,
  output        hitLD_0,
  output        missLD_0,
  output        _T_294_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
`endif // RANDOMIZE_REG_INIT
  wire  cache_clock; // @[programmableCache.scala 52:26]
  wire  cache_reset; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_0_req_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_cpu_0_req_bits_addr; // @[programmableCache.scala 52:26]
  wire [63:0] cache_io_cpu_0_req_bits_data; // @[programmableCache.scala 52:26]
  wire [27:0] cache_io_cpu_0_req_bits_command; // @[programmableCache.scala 52:26]
  wire [2:0] cache_io_cpu_0_req_bits_way; // @[programmableCache.scala 52:26]
  wire [2:0] cache_io_cpu_0_req_bits_replaceWay; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_0_resp_valid; // @[programmableCache.scala 52:26]
  wire  cache_io_cpu_0_resp_bits_iswrite; // @[programmableCache.scala 52:26]
  wire [2:0] cache_io_cpu_0_resp_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_probe_req_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_probe_req_bits_addr; // @[programmableCache.scala 52:26]
  wire [27:0] cache_io_probe_req_bits_command; // @[programmableCache.scala 52:26]
  wire  cache_io_probe_resp_valid; // @[programmableCache.scala 52:26]
  wire [2:0] cache_io_probe_resp_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_probe_multiWay_valid; // @[programmableCache.scala 52:26]
  wire [2:0] cache_io_probe_multiWay_bits_way_0; // @[programmableCache.scala 52:26]
  wire [2:0] cache_io_probe_multiWay_bits_way_1; // @[programmableCache.scala 52:26]
  wire [2:0] cache_io_probe_multiWay_bits_way_2; // @[programmableCache.scala 52:26]
  wire [2:0] cache_io_probe_multiWay_bits_way_3; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_probe_multiWay_bits_addr; // @[programmableCache.scala 52:26]
  wire  cache_io_bipassLD_in_valid; // @[programmableCache.scala 52:26]
  wire [31:0] cache_io_bipassLD_in_bits_addr; // @[programmableCache.scala 52:26]
  wire [3:0] cache_io_bipassLD_in_bits_way; // @[programmableCache.scala 52:26]
  wire  cache_io_bipassLD_out_valid; // @[programmableCache.scala 52:26]
  wire [63:0] cache_io_bipassLD_out_bits_data; // @[programmableCache.scala 52:26]
  wire  tbe_clock; // @[programmableCache.scala 53:26]
  wire  tbe_reset; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_0_valid; // @[programmableCache.scala 53:26]
  wire [63:0] tbe_io_write_0_bits_addr; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_0_bits_command; // @[programmableCache.scala 53:26]
  wire  tbe_io_write_0_bits_mask; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_write_0_bits_inputTBE_state_state; // @[programmableCache.scala 53:26]
  wire [3:0] tbe_io_write_0_bits_inputTBE_way; // @[programmableCache.scala 53:26]
  wire [31:0] tbe_io_write_0_bits_inputTBE_fields_0; // @[programmableCache.scala 53:26]
  wire  tbe_io_read_valid; // @[programmableCache.scala 53:26]
  wire [63:0] tbe_io_read_bits_addr; // @[programmableCache.scala 53:26]
  wire [1:0] tbe_io_outputTBE_bits_state_state; // @[programmableCache.scala 53:26]
  wire [3:0] tbe_io_outputTBE_bits_way; // @[programmableCache.scala 53:26]
  wire [31:0] tbe_io_outputTBE_bits_fields_0; // @[programmableCache.scala 53:26]
  wire  tbe_io_isFull; // @[programmableCache.scala 53:26]
  wire  lockMem_clock; // @[programmableCache.scala 54:26]
  wire  lockMem_reset; // @[programmableCache.scala 54:26]
  wire  lockMem_io_lock_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_lock_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  lockMem_io_probe_out_valid; // @[programmableCache.scala 54:26]
  wire  lockMem_io_probe_out_bits; // @[programmableCache.scala 54:26]
  wire  lockMem_io_probe_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_probe_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  lockMem_io_unLock_0_in_valid; // @[programmableCache.scala 54:26]
  wire [31:0] lockMem_io_unLock_0_in_bits_addr; // @[programmableCache.scala 54:26]
  wire  stateMem_clock; // @[programmableCache.scala 55:27]
  wire  stateMem_reset; // @[programmableCache.scala 55:27]
  wire  stateMem_io_in_0_valid; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_in_0_bits_state_state; // @[programmableCache.scala 55:27]
  wire [31:0] stateMem_io_in_0_bits_addr; // @[programmableCache.scala 55:27]
  wire [2:0] stateMem_io_in_0_bits_way; // @[programmableCache.scala 55:27]
  wire  stateMem_io_in_1_valid; // @[programmableCache.scala 55:27]
  wire [31:0] stateMem_io_in_1_bits_addr; // @[programmableCache.scala 55:27]
  wire [2:0] stateMem_io_in_1_bits_way; // @[programmableCache.scala 55:27]
  wire  stateMem_io_out_valid; // @[programmableCache.scala 55:27]
  wire [1:0] stateMem_io_out_bits_state; // @[programmableCache.scala 55:27]
  wire  pc_clock; // @[programmableCache.scala 56:26]
  wire  pc_reset; // @[programmableCache.scala 56:26]
  wire  pc_io_write_ready; // @[programmableCache.scala 56:26]
  wire  pc_io_write_valid; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_write_bits_addr; // @[programmableCache.scala 56:26]
  wire [2:0] pc_io_write_bits_way; // @[programmableCache.scala 56:26]
  wire [63:0] pc_io_write_bits_data; // @[programmableCache.scala 56:26]
  wire [2:0] pc_io_write_bits_replaceWay; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_write_bits_tbeFields_0; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_write_bits_pc; // @[programmableCache.scala 56:26]
  wire [2:0] pc_io_read_0_in_bits_data_way; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_0_in_bits_data_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_0_in_bits_data_valid; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_0_out_bits_addr; // @[programmableCache.scala 56:26]
  wire [2:0] pc_io_read_0_out_bits_way; // @[programmableCache.scala 56:26]
  wire [63:0] pc_io_read_0_out_bits_data; // @[programmableCache.scala 56:26]
  wire [2:0] pc_io_read_0_out_bits_replaceWay; // @[programmableCache.scala 56:26]
  wire [31:0] pc_io_read_0_out_bits_tbeFields_0; // @[programmableCache.scala 56:26]
  wire [15:0] pc_io_read_0_out_bits_pc; // @[programmableCache.scala 56:26]
  wire  pc_io_read_0_out_bits_valid; // @[programmableCache.scala 56:26]
  wire  pc_io_isFull; // @[programmableCache.scala 56:26]
  wire  inputArbiter_io_in_0_valid; // @[programmableCache.scala 57:33]
  wire [1:0] inputArbiter_io_in_0_bits_event; // @[programmableCache.scala 57:33]
  wire [31:0] inputArbiter_io_in_0_bits_addr; // @[programmableCache.scala 57:33]
  wire [63:0] inputArbiter_io_in_0_bits_data; // @[programmableCache.scala 57:33]
  wire  inputArbiter_io_in_1_ready; // @[programmableCache.scala 57:33]
  wire  inputArbiter_io_in_1_valid; // @[programmableCache.scala 57:33]
  wire [1:0] inputArbiter_io_in_1_bits_event; // @[programmableCache.scala 57:33]
  wire [31:0] inputArbiter_io_in_1_bits_addr; // @[programmableCache.scala 57:33]
  wire [63:0] inputArbiter_io_in_1_bits_data; // @[programmableCache.scala 57:33]
  wire  inputArbiter_io_in_2_valid; // @[programmableCache.scala 57:33]
  wire [1:0] inputArbiter_io_in_2_bits_event; // @[programmableCache.scala 57:33]
  wire [31:0] inputArbiter_io_in_2_bits_addr; // @[programmableCache.scala 57:33]
  wire [63:0] inputArbiter_io_in_2_bits_data; // @[programmableCache.scala 57:33]
  wire  inputArbiter_io_in_3_valid; // @[programmableCache.scala 57:33]
  wire [1:0] inputArbiter_io_in_3_bits_event; // @[programmableCache.scala 57:33]
  wire [31:0] inputArbiter_io_in_3_bits_addr; // @[programmableCache.scala 57:33]
  wire [63:0] inputArbiter_io_in_3_bits_data; // @[programmableCache.scala 57:33]
  wire  inputArbiter_io_out_ready; // @[programmableCache.scala 57:33]
  wire  inputArbiter_io_out_valid; // @[programmableCache.scala 57:33]
  wire [1:0] inputArbiter_io_out_bits_event; // @[programmableCache.scala 57:33]
  wire [31:0] inputArbiter_io_out_bits_addr; // @[programmableCache.scala 57:33]
  wire [63:0] inputArbiter_io_out_bits_data; // @[programmableCache.scala 57:33]
  wire [1:0] inputArbiter_io_chosen; // @[programmableCache.scala 57:33]
  wire  outReqArbiter_io_in_0_valid; // @[programmableCache.scala 58:33]
  wire [31:0] outReqArbiter_io_in_0_bits_req_addr; // @[programmableCache.scala 58:33]
  wire [7:0] outReqArbiter_io_in_0_bits_req_inst; // @[programmableCache.scala 58:33]
  wire [63:0] outReqArbiter_io_in_0_bits_req_data; // @[programmableCache.scala 58:33]
  wire  outReqArbiter_io_out_valid; // @[programmableCache.scala 58:33]
  wire [31:0] outReqArbiter_io_out_bits_req_addr; // @[programmableCache.scala 58:33]
  wire [7:0] outReqArbiter_io_out_bits_req_inst; // @[programmableCache.scala 58:33]
  wire [63:0] outReqArbiter_io_out_bits_req_data; // @[programmableCache.scala 58:33]
  wire  outRespArbiter_io_in_0_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_in_0_bits_addr; // @[programmableCache.scala 59:33]
  wire  outRespArbiter_io_in_1_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_in_1_bits_addr; // @[programmableCache.scala 59:33]
  wire  outRespArbiter_io_out_valid; // @[programmableCache.scala 59:33]
  wire [31:0] outRespArbiter_io_out_bits_addr; // @[programmableCache.scala 59:33]
  wire  feedbackArbiter_io_in_0_ready; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_in_0_valid; // @[programmableCache.scala 60:34]
  wire [1:0] feedbackArbiter_io_in_0_bits_event; // @[programmableCache.scala 60:34]
  wire [31:0] feedbackArbiter_io_in_0_bits_addr; // @[programmableCache.scala 60:34]
  wire [63:0] feedbackArbiter_io_in_0_bits_data; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_out_ready; // @[programmableCache.scala 60:34]
  wire  feedbackArbiter_io_out_valid; // @[programmableCache.scala 60:34]
  wire [1:0] feedbackArbiter_io_out_bits_event; // @[programmableCache.scala 60:34]
  wire [31:0] feedbackArbiter_io_out_bits_addr; // @[programmableCache.scala 60:34]
  wire [63:0] feedbackArbiter_io_out_bits_data; // @[programmableCache.scala 60:34]
  wire  input__clock; // @[programmableCache.scala 90:23]
  wire  input__reset; // @[programmableCache.scala 90:23]
  wire  input__io_enq_ready; // @[programmableCache.scala 90:23]
  wire  input__io_enq_valid; // @[programmableCache.scala 90:23]
  wire [1:0] input__io_enq_bits_inst_event; // @[programmableCache.scala 90:23]
  wire [31:0] input__io_enq_bits_inst_addr; // @[programmableCache.scala 90:23]
  wire [63:0] input__io_enq_bits_inst_data; // @[programmableCache.scala 90:23]
  wire [1:0] input__io_enq_bits_tbeOut_state_state; // @[programmableCache.scala 90:23]
  wire [3:0] input__io_enq_bits_tbeOut_way; // @[programmableCache.scala 90:23]
  wire [31:0] input__io_enq_bits_tbeOut_fields_0; // @[programmableCache.scala 90:23]
  wire  input__io_deq_ready; // @[programmableCache.scala 90:23]
  wire  input__io_deq_valid; // @[programmableCache.scala 90:23]
  wire [1:0] input__io_deq_bits_inst_event; // @[programmableCache.scala 90:23]
  wire [31:0] input__io_deq_bits_inst_addr; // @[programmableCache.scala 90:23]
  wire [63:0] input__io_deq_bits_inst_data; // @[programmableCache.scala 90:23]
  wire [1:0] input__io_deq_bits_tbeOut_state_state; // @[programmableCache.scala 90:23]
  wire [3:0] input__io_deq_bits_tbeOut_way; // @[programmableCache.scala 90:23]
  wire [31:0] input__io_deq_bits_tbeOut_fields_0; // @[programmableCache.scala 90:23]
  wire  respPortQueue_0_clock; // @[programmableCache.scala 93:27]
  wire  respPortQueue_0_reset; // @[programmableCache.scala 93:27]
  wire  respPortQueue_0_io_enq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_0_io_enq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_0_io_enq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_0_io_enq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_0_io_enq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_0_io_deq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_0_io_deq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_0_io_deq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_0_io_deq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_0_io_deq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_1_clock; // @[programmableCache.scala 93:27]
  wire  respPortQueue_1_reset; // @[programmableCache.scala 93:27]
  wire  respPortQueue_1_io_enq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_1_io_enq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_1_io_enq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_1_io_enq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_1_io_enq_bits_data; // @[programmableCache.scala 93:27]
  wire  respPortQueue_1_io_deq_ready; // @[programmableCache.scala 93:27]
  wire  respPortQueue_1_io_deq_valid; // @[programmableCache.scala 93:27]
  wire [1:0] respPortQueue_1_io_deq_bits_event; // @[programmableCache.scala 93:27]
  wire [31:0] respPortQueue_1_io_deq_bits_addr; // @[programmableCache.scala 93:27]
  wire [63:0] respPortQueue_1_io_deq_bits_data; // @[programmableCache.scala 93:27]
  wire  reqPortQueue_0_clock; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_0_reset; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_0_io_enq_ready; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_0_io_enq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_0_io_enq_bits_addr; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_0_io_enq_bits_data; // @[programmableCache.scala 98:27]
  wire  reqPortQueue_0_io_deq_valid; // @[programmableCache.scala 98:27]
  wire [31:0] reqPortQueue_0_io_deq_bits_addr; // @[programmableCache.scala 98:27]
  wire [7:0] reqPortQueue_0_io_deq_bits_inst; // @[programmableCache.scala 98:27]
  wire [63:0] reqPortQueue_0_io_deq_bits_data; // @[programmableCache.scala 98:27]
  wire  feedbackInQueue_0_clock; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_0_reset; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_0_io_enq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_0_io_enq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_0_io_enq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_0_io_enq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_0_io_enq_bits_data; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_0_io_deq_ready; // @[programmableCache.scala 104:27]
  wire  feedbackInQueue_0_io_deq_valid; // @[programmableCache.scala 104:27]
  wire [1:0] feedbackInQueue_0_io_deq_bits_event; // @[programmableCache.scala 104:27]
  wire [31:0] feedbackInQueue_0_io_deq_bits_addr; // @[programmableCache.scala 104:27]
  wire [63:0] feedbackInQueue_0_io_deq_bits_data; // @[programmableCache.scala 104:27]
  wire  probeWay_clock; // @[programmableCache.scala 108:26]
  wire  probeWay_reset; // @[programmableCache.scala 108:26]
  wire  probeWay_io_enq_ready; // @[programmableCache.scala 108:26]
  wire  probeWay_io_enq_valid; // @[programmableCache.scala 108:26]
  wire [2:0] probeWay_io_enq_bits; // @[programmableCache.scala 108:26]
  wire  probeWay_io_deq_ready; // @[programmableCache.scala 108:26]
  wire  probeWay_io_deq_valid; // @[programmableCache.scala 108:26]
  wire [2:0] probeWay_io_deq_bits; // @[programmableCache.scala 108:26]
  wire  feedbackOutQueue_clock; // @[programmableCache.scala 165:34]
  wire  feedbackOutQueue_reset; // @[programmableCache.scala 165:34]
  wire  feedbackOutQueue_io_enq_ready; // @[programmableCache.scala 165:34]
  wire  feedbackOutQueue_io_enq_valid; // @[programmableCache.scala 165:34]
  wire [1:0] feedbackOutQueue_io_enq_bits_event; // @[programmableCache.scala 165:34]
  wire [31:0] feedbackOutQueue_io_enq_bits_addr; // @[programmableCache.scala 165:34]
  wire [63:0] feedbackOutQueue_io_enq_bits_data; // @[programmableCache.scala 165:34]
  wire  feedbackOutQueue_io_deq_ready; // @[programmableCache.scala 165:34]
  wire  feedbackOutQueue_io_deq_valid; // @[programmableCache.scala 165:34]
  wire [1:0] feedbackOutQueue_io_deq_bits_event; // @[programmableCache.scala 165:34]
  wire [31:0] feedbackOutQueue_io_deq_bits_addr; // @[programmableCache.scala 165:34]
  wire [63:0] feedbackOutQueue_io_deq_bits_data; // @[programmableCache.scala 165:34]
  wire  routineQueue_clock; // @[programmableCache.scala 166:30]
  wire  routineQueue_reset; // @[programmableCache.scala 166:30]
  wire  routineQueue_io_enq_ready; // @[programmableCache.scala 166:30]
  wire  routineQueue_io_enq_valid; // @[programmableCache.scala 166:30]
  wire [15:0] routineQueue_io_enq_bits; // @[programmableCache.scala 166:30]
  wire  routineQueue_io_deq_ready; // @[programmableCache.scala 166:30]
  wire  routineQueue_io_deq_valid; // @[programmableCache.scala 166:30]
  wire [15:0] routineQueue_io_deq_bits; // @[programmableCache.scala 166:30]
  wire  actionReg_0_clock; // @[programmableCache.scala 169:32]
  wire  actionReg_0_reset; // @[programmableCache.scala 169:32]
  wire  actionReg_0_io_enq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_0_io_enq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_0_io_enq_bits_addr; // @[programmableCache.scala 169:32]
  wire [2:0] actionReg_0_io_enq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_0_io_enq_bits_data; // @[programmableCache.scala 169:32]
  wire [2:0] actionReg_0_io_enq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_0_io_enq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_0_io_enq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_0_io_enq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  actionReg_0_io_deq_ready; // @[programmableCache.scala 169:32]
  wire  actionReg_0_io_deq_valid; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_0_io_deq_bits_addr; // @[programmableCache.scala 169:32]
  wire [2:0] actionReg_0_io_deq_bits_way; // @[programmableCache.scala 169:32]
  wire [63:0] actionReg_0_io_deq_bits_data; // @[programmableCache.scala 169:32]
  wire [2:0] actionReg_0_io_deq_bits_replaceWay; // @[programmableCache.scala 169:32]
  wire [31:0] actionReg_0_io_deq_bits_tbeFields_0; // @[programmableCache.scala 169:32]
  wire [27:0] actionReg_0_io_deq_bits_action_signals; // @[programmableCache.scala 169:32]
  wire [3:0] actionReg_0_io_deq_bits_action_actionType; // @[programmableCache.scala 169:32]
  wire  mimoQ_clock; // @[programmableCache.scala 173:24]
  wire  mimoQ_reset; // @[programmableCache.scala 173:24]
  wire  mimoQ_io_enq_ready; // @[programmableCache.scala 173:24]
  wire  mimoQ_io_enq_valid; // @[programmableCache.scala 173:24]
  wire [2:0] mimoQ_io_enq_bits_0_way; // @[programmableCache.scala 173:24]
  wire [31:0] mimoQ_io_enq_bits_0_addr; // @[programmableCache.scala 173:24]
  wire [2:0] mimoQ_io_enq_bits_1_way; // @[programmableCache.scala 173:24]
  wire [31:0] mimoQ_io_enq_bits_1_addr; // @[programmableCache.scala 173:24]
  wire [2:0] mimoQ_io_enq_bits_2_way; // @[programmableCache.scala 173:24]
  wire [31:0] mimoQ_io_enq_bits_2_addr; // @[programmableCache.scala 173:24]
  wire [2:0] mimoQ_io_enq_bits_3_way; // @[programmableCache.scala 173:24]
  wire [31:0] mimoQ_io_enq_bits_3_addr; // @[programmableCache.scala 173:24]
  wire  mimoQ_io_deq_valid; // @[programmableCache.scala 173:24]
  wire [2:0] mimoQ_io_deq_bits_0_way; // @[programmableCache.scala 173:24]
  wire [31:0] mimoQ_io_deq_bits_0_addr; // @[programmableCache.scala 173:24]
  wire [7:0] mimoQ_io_count; // @[programmableCache.scala 173:24]
  wire  compUnit_0_clock; // @[programmableCache.scala 177:27]
  wire  compUnit_0_reset; // @[programmableCache.scala 177:27]
  wire  compUnit_0_io_instruction_valid; // @[programmableCache.scala 177:27]
  wire [27:0] compUnit_0_io_instruction_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_0_io_clear; // @[programmableCache.scala 177:27]
  wire  compUnit_0_io_op1_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_0_io_op1_bits; // @[programmableCache.scala 177:27]
  wire  compUnit_0_io_op2_valid; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_0_io_op2_bits; // @[programmableCache.scala 177:27]
  wire [15:0] compUnit_0_io_pc; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_0_io_reg_file_0; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_0_io_reg_file_1; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_0_io_reg_file_2; // @[programmableCache.scala 177:27]
  wire [63:0] compUnit_0_io_reg_file_3; // @[programmableCache.scala 177:27]
  wire [63:0] compUnitInput1_0_io_in_hardCoded; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_0_io_in_data; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_0_io_in_tbe; // @[programmableCache.scala 182:30]
  wire [1:0] compUnitInput1_0_io_in_select; // @[programmableCache.scala 182:30]
  wire  compUnitInput1_0_io_out_valid; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput1_0_io_out_bits; // @[programmableCache.scala 182:30]
  wire [63:0] compUnitInput2_0_io_in_hardCoded; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_0_io_in_data; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_0_io_in_tbe; // @[programmableCache.scala 188:30]
  wire [1:0] compUnitInput2_0_io_in_select; // @[programmableCache.scala 188:30]
  wire  compUnitInput2_0_io_out_valid; // @[programmableCache.scala 188:30]
  wire [63:0] compUnitInput2_0_io_out_bits; // @[programmableCache.scala 188:30]
  wire  _T_95 = input__io_deq_bits_tbeOut_state_state != 2'h0; // @[programmableCache.scala 293:55]
  wire [1:0] _T_96 = stateMem_io_out_valid ? stateMem_io_out_bits_state : 2'h0; // @[programmableCache.scala 293:120]
  wire [1:0] state = _T_95 ? input__io_deq_bits_tbeOut_state_state : _T_96; // @[programmableCache.scala 293:17]
  wire [3:0] routine = {input__io_deq_bits_inst_event,state}; // @[Cat.scala 29:58]
  reg  instUsed; // @[programmableCache.scala 197:27]
  reg [5:0] replStateReg_0; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_1; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_2; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_3; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_4; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_5; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_6; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_7; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_8; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_9; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_10; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_11; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_12; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_13; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_14; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_15; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_16; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_17; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_18; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_19; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_20; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_21; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_22; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_23; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_24; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_25; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_26; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_27; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_28; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_29; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_30; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_31; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_32; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_33; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_34; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_35; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_36; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_37; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_38; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_39; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_40; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_41; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_42; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_43; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_44; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_45; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_46; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_47; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_48; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_49; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_50; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_51; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_52; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_53; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_54; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_55; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_56; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_57; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_58; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_59; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_60; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_61; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_62; // @[programmableCache.scala 204:31]
  reg [5:0] replStateReg_63; // @[programmableCache.scala 204:31]
  wire [31:0] _GEN_385 = {{24'd0}, actionReg_0_io_deq_bits_action_signals[7:0]}; // @[programmableCache.scala 247:78]
  wire [63:0] _GEN_386 = {{60'd0}, actionReg_0_io_deq_bits_action_signals[11:8]}; // @[programmableCache.scala 249:78]
  wire  isLocked = lockMem_io_probe_out_valid & lockMem_io_probe_out_bits; // @[programmableCache.scala 323:21]
  wire  stallInput = isLocked | tbe_io_isFull; // @[programmableCache.scala 260:28]
  wire  _T_47 = 2'h1 == input__io_deq_bits_inst_event; // @[programmableCache.scala 264:35]
  wire  _T_48 = 2'h0 == input__io_deq_bits_inst_event; // @[programmableCache.scala 264:35]
  wire  hitEvent = _T_47 | _T_48; // @[programmableCache.scala 264:35]
  wire  _T_84 = ~tbe_io_isFull; // @[programmableCache.scala 284:48]
  wire  _T_85 = input__io_enq_ready & _T_84; // @[programmableCache.scala 284:45]
  wire  _T_86 = ~stallInput; // @[programmableCache.scala 284:66]
  wire  instruction_ready = _T_85 & _T_86; // @[programmableCache.scala 284:63]
  wire  instruction_valid = inputArbiter_io_out_valid; // @[programmableCache.scala 110:27 programmableCache.scala 252:17]
  wire  _T_52 = instruction_ready & instruction_valid; // @[Decoupled.scala 40:37]
  wire [1:0] instruction_bits_event = inputArbiter_io_out_bits_event; // @[programmableCache.scala 110:27 programmableCache.scala 252:17]
  wire  _T_53 = 2'h1 == instruction_bits_event; // @[programmableCache.scala 267:59]
  wire  _T_54 = 2'h0 == instruction_bits_event; // @[programmableCache.scala 267:59]
  wire  _T_56 = _T_53 | _T_54; // @[programmableCache.scala 267:59]
  wire  probeStart = _T_52 & _T_56; // @[programmableCache.scala 267:38]
  wire  getState = input__io_deq_ready & input__io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_62 = probeWay_io_deq_bits != 3'h4; // @[programmableCache.scala 275:46]
  wire  _T_63 = getState & _T_62; // @[programmableCache.scala 275:21]
  wire  _T_64 = stateMem_io_out_bits_state == 2'h2; // @[programmableCache.scala 275:90]
  wire  hit = _T_63 & _T_64; // @[programmableCache.scala 275:59]
  wire  _T_66 = hit & hitEvent; // @[programmableCache.scala 276:20]
  wire  _T_67 = getState & hitEvent; // @[programmableCache.scala 277:24]
  wire  _T_68 = stateMem_io_out_bits_state == 2'h0; // @[programmableCache.scala 277:71]
  wire  _T_69 = _T_67 & _T_68; // @[programmableCache.scala 277:39]
  wire  _T_71 = inputArbiter_io_chosen == 2'h0; // @[programmableCache.scala 279:77]
  wire  _T_72 = _T_52 & _T_71; // @[programmableCache.scala 279:51]
  wire  _T_74 = inputArbiter_io_chosen == 2'h3; // @[programmableCache.scala 280:76]
  wire  _T_75 = _T_52 & _T_74; // @[programmableCache.scala 280:50]
  wire  _T_77 = inputArbiter_io_chosen == 2'h2; // @[programmableCache.scala 281:77]
  wire  _T_80 = ~_T_52; // @[programmableCache.scala 283:20]
  wire  _T_81 = input__io_enq_ready & input__io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_82 = _T_81 | instUsed; // @[programmableCache.scala 283:63]
  wire  _T_83 = _T_80 & _T_82; // @[programmableCache.scala 283:40]
  wire  _T_88 = ~instUsed; // @[programmableCache.scala 286:48]
  wire  _T_89 = instruction_valid & _T_88; // @[programmableCache.scala 286:45]
  wire  _T_91 = _T_89 & _T_84; // @[programmableCache.scala 286:58]
  wire  maskField_0 = actionReg_0_io_deq_bits_action_signals[2]; // @[Gem5CacheLogic.scala 114:54]
  wire  _T_98 = ~maskField_0; // @[programmableCache.scala 303:84]
  wire [63:0] _GEN_377 = compUnit_0_io_reg_file_0; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_378 = 2'h1 == actionReg_0_io_deq_bits_action_signals[4:3] ? compUnit_0_io_reg_file_1 : _GEN_377; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_379 = 2'h2 == actionReg_0_io_deq_bits_action_signals[4:3] ? compUnit_0_io_reg_file_2 : _GEN_378; // @[programmableCache.scala 417:31]
  wire [63:0] _GEN_380 = 2'h3 == actionReg_0_io_deq_bits_action_signals[4:3] ? compUnit_0_io_reg_file_3 : _GEN_379; // @[programmableCache.scala 417:31]
  wire [31:0] tbeFieldUpdateSrc_0 = _GEN_380[31:0]; // @[programmableCache.scala 138:33 programmableCache.scala 417:31]
  wire  _T_204 = actionReg_0_io_deq_bits_action_actionType == 4'h3; // @[programmableCache.scala 373:73]
  wire  isStateAction_0 = _T_204 & actionReg_0_io_deq_valid; // @[programmableCache.scala 373:82]
  wire [1:0] tbeAction_0 = actionReg_0_io_deq_bits_action_signals[1:0]; // @[Gem5CacheLogic.scala 115:54]
  wire  _T_198 = actionReg_0_io_deq_bits_action_actionType == 4'h1; // @[programmableCache.scala 370:73]
  wire  isTBEAction_0 = _T_198 & actionReg_0_io_deq_valid; // @[programmableCache.scala 370:82]
  wire [4:0] _GEN_1 = 4'h1 == routine ? 5'h0 : 5'h1; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_2 = 4'h2 == routine ? 5'h1a : _GEN_1; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_3 = 4'h3 == routine ? 5'h0 : _GEN_2; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_4 = 4'h4 == routine ? 5'h8 : _GEN_3; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_5 = 4'h5 == routine ? 5'h0 : _GEN_4; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_6 = 4'h6 == routine ? 5'h0 : _GEN_5; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_7 = 4'h7 == routine ? 5'h0 : _GEN_6; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_8 = 4'h8 == routine ? 5'h1d : _GEN_7; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_9 = 4'h9 == routine ? 5'h11 : _GEN_8; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_10 = 4'ha == routine ? 5'h0 : _GEN_9; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_11 = 4'hb == routine ? 5'h0 : _GEN_10; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_12 = 4'hc == routine ? 5'h16 : _GEN_11; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_13 = 4'hd == routine ? 5'h0 : _GEN_12; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_14 = 4'he == routine ? 5'h0 : _GEN_13; // @[programmableCache.scala 349:30]
  wire [4:0] _GEN_15 = 4'hf == routine ? 5'h0 : _GEN_14; // @[programmableCache.scala 349:30]
  wire [31:0] addrReplacer = {{26'd0}, input__io_deq_bits_inst_addr[8:3]}; // @[programmableCache.scala 207:28 programmableCache.scala 356:18]
  wire [5:0] _GEN_17 = 6'h1 == addrReplacer[5:0] ? replStateReg_1 : replStateReg_0; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_18 = 6'h2 == addrReplacer[5:0] ? replStateReg_2 : _GEN_17; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_19 = 6'h3 == addrReplacer[5:0] ? replStateReg_3 : _GEN_18; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_20 = 6'h4 == addrReplacer[5:0] ? replStateReg_4 : _GEN_19; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_21 = 6'h5 == addrReplacer[5:0] ? replStateReg_5 : _GEN_20; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_22 = 6'h6 == addrReplacer[5:0] ? replStateReg_6 : _GEN_21; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_23 = 6'h7 == addrReplacer[5:0] ? replStateReg_7 : _GEN_22; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_24 = 6'h8 == addrReplacer[5:0] ? replStateReg_8 : _GEN_23; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_25 = 6'h9 == addrReplacer[5:0] ? replStateReg_9 : _GEN_24; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_26 = 6'ha == addrReplacer[5:0] ? replStateReg_10 : _GEN_25; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_27 = 6'hb == addrReplacer[5:0] ? replStateReg_11 : _GEN_26; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_28 = 6'hc == addrReplacer[5:0] ? replStateReg_12 : _GEN_27; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_29 = 6'hd == addrReplacer[5:0] ? replStateReg_13 : _GEN_28; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_30 = 6'he == addrReplacer[5:0] ? replStateReg_14 : _GEN_29; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_31 = 6'hf == addrReplacer[5:0] ? replStateReg_15 : _GEN_30; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_32 = 6'h10 == addrReplacer[5:0] ? replStateReg_16 : _GEN_31; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_33 = 6'h11 == addrReplacer[5:0] ? replStateReg_17 : _GEN_32; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_34 = 6'h12 == addrReplacer[5:0] ? replStateReg_18 : _GEN_33; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_35 = 6'h13 == addrReplacer[5:0] ? replStateReg_19 : _GEN_34; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_36 = 6'h14 == addrReplacer[5:0] ? replStateReg_20 : _GEN_35; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_37 = 6'h15 == addrReplacer[5:0] ? replStateReg_21 : _GEN_36; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_38 = 6'h16 == addrReplacer[5:0] ? replStateReg_22 : _GEN_37; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_39 = 6'h17 == addrReplacer[5:0] ? replStateReg_23 : _GEN_38; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_40 = 6'h18 == addrReplacer[5:0] ? replStateReg_24 : _GEN_39; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_41 = 6'h19 == addrReplacer[5:0] ? replStateReg_25 : _GEN_40; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_42 = 6'h1a == addrReplacer[5:0] ? replStateReg_26 : _GEN_41; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_43 = 6'h1b == addrReplacer[5:0] ? replStateReg_27 : _GEN_42; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_44 = 6'h1c == addrReplacer[5:0] ? replStateReg_28 : _GEN_43; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_45 = 6'h1d == addrReplacer[5:0] ? replStateReg_29 : _GEN_44; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_46 = 6'h1e == addrReplacer[5:0] ? replStateReg_30 : _GEN_45; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_47 = 6'h1f == addrReplacer[5:0] ? replStateReg_31 : _GEN_46; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_48 = 6'h20 == addrReplacer[5:0] ? replStateReg_32 : _GEN_47; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_49 = 6'h21 == addrReplacer[5:0] ? replStateReg_33 : _GEN_48; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_50 = 6'h22 == addrReplacer[5:0] ? replStateReg_34 : _GEN_49; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_51 = 6'h23 == addrReplacer[5:0] ? replStateReg_35 : _GEN_50; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_52 = 6'h24 == addrReplacer[5:0] ? replStateReg_36 : _GEN_51; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_53 = 6'h25 == addrReplacer[5:0] ? replStateReg_37 : _GEN_52; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_54 = 6'h26 == addrReplacer[5:0] ? replStateReg_38 : _GEN_53; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_55 = 6'h27 == addrReplacer[5:0] ? replStateReg_39 : _GEN_54; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_56 = 6'h28 == addrReplacer[5:0] ? replStateReg_40 : _GEN_55; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_57 = 6'h29 == addrReplacer[5:0] ? replStateReg_41 : _GEN_56; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_58 = 6'h2a == addrReplacer[5:0] ? replStateReg_42 : _GEN_57; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_59 = 6'h2b == addrReplacer[5:0] ? replStateReg_43 : _GEN_58; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_60 = 6'h2c == addrReplacer[5:0] ? replStateReg_44 : _GEN_59; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_61 = 6'h2d == addrReplacer[5:0] ? replStateReg_45 : _GEN_60; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_62 = 6'h2e == addrReplacer[5:0] ? replStateReg_46 : _GEN_61; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_63 = 6'h2f == addrReplacer[5:0] ? replStateReg_47 : _GEN_62; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_64 = 6'h30 == addrReplacer[5:0] ? replStateReg_48 : _GEN_63; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_65 = 6'h31 == addrReplacer[5:0] ? replStateReg_49 : _GEN_64; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_66 = 6'h32 == addrReplacer[5:0] ? replStateReg_50 : _GEN_65; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_67 = 6'h33 == addrReplacer[5:0] ? replStateReg_51 : _GEN_66; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_68 = 6'h34 == addrReplacer[5:0] ? replStateReg_52 : _GEN_67; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_69 = 6'h35 == addrReplacer[5:0] ? replStateReg_53 : _GEN_68; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_70 = 6'h36 == addrReplacer[5:0] ? replStateReg_54 : _GEN_69; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_71 = 6'h37 == addrReplacer[5:0] ? replStateReg_55 : _GEN_70; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_72 = 6'h38 == addrReplacer[5:0] ? replStateReg_56 : _GEN_71; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_73 = 6'h39 == addrReplacer[5:0] ? replStateReg_57 : _GEN_72; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_74 = 6'h3a == addrReplacer[5:0] ? replStateReg_58 : _GEN_73; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_75 = 6'h3b == addrReplacer[5:0] ? replStateReg_59 : _GEN_74; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_76 = 6'h3c == addrReplacer[5:0] ? replStateReg_60 : _GEN_75; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_77 = 6'h3d == addrReplacer[5:0] ? replStateReg_61 : _GEN_76; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_78 = 6'h3e == addrReplacer[5:0] ? replStateReg_62 : _GEN_77; // @[Replacement.scala 97:41]
  wire [5:0] _GEN_79 = 6'h3f == addrReplacer[5:0] ? replStateReg_63 : _GEN_78; // @[Replacement.scala 97:41]
  wire [3:0] _T_112 = {_GEN_79[2:0],1'h0}; // @[Cat.scala 29:58]
  wire [3:0] _T_114 = {_GEN_79[4:3],2'h0}; // @[Cat.scala 29:58]
  wire [3:0] _T_116 = {_GEN_79[5],3'h0}; // @[Cat.scala 29:58]
  wire  _T_118 = &_T_112[3:1]; // @[Replacement.scala 133:103]
  wire  _T_121 = &_T_114[3:2]; // @[Replacement.scala 133:103]
  wire  _T_123 = ~_T_112[1]; // @[Replacement.scala 134:89]
  wire  _T_125 = ~_T_114[1]; // @[Replacement.scala 134:89]
  wire  _T_127 = ~_T_116[1]; // @[Replacement.scala 134:89]
  wire  _T_128 = _T_123 & _T_125; // @[Replacement.scala 134:105]
  wire  _T_129 = _T_128 & _T_127; // @[Replacement.scala 134:105]
  wire  _T_130 = _T_121 & _T_129; // @[Replacement.scala 135:28]
  wire  _T_132 = &_T_116[3]; // @[Replacement.scala 133:103]
  wire  _T_134 = ~_T_112[2]; // @[Replacement.scala 134:89]
  wire  _T_136 = ~_T_114[2]; // @[Replacement.scala 134:89]
  wire  _T_138 = ~_T_116[2]; // @[Replacement.scala 134:89]
  wire  _T_139 = _T_134 & _T_136; // @[Replacement.scala 134:105]
  wire  _T_140 = _T_139 & _T_138; // @[Replacement.scala 134:105]
  wire  _T_141 = _T_132 & _T_140; // @[Replacement.scala 135:28]
  wire  _T_143 = ~_T_112[3]; // @[Replacement.scala 134:89]
  wire  _T_145 = ~_T_114[3]; // @[Replacement.scala 134:89]
  wire  _T_147 = ~_T_116[3]; // @[Replacement.scala 134:89]
  wire  _T_148 = _T_143 & _T_145; // @[Replacement.scala 134:105]
  wire  _T_149 = _T_148 & _T_147; // @[Replacement.scala 134:105]
  wire [3:0] _T_153 = {_T_149,_T_141,_T_130,_T_118}; // @[Cat.scala 29:58]
  wire  _T_156 = |_T_153[3:2]; // @[OneHot.scala 32:14]
  wire [1:0] _T_157 = _T_153[3:2] | _T_153[1:0]; // @[OneHot.scala 32:28]
  wire [1:0] _T_159 = {_T_156,_T_157[1]}; // @[Cat.scala 29:58]
  wire [5:0] replacerWayWire = {{4'd0}, _T_159}; // @[programmableCache.scala 205:31 programmableCache.scala 357:21]
  wire [3:0] _T_171 = 4'h1 << replacerWayWire[1:0]; // @[OneHot.scala 65:12]
  wire  _T_173 = 6'h0 == replacerWayWire; // @[Replacement.scala 111:25]
  wire [3:0] _T_174 = _T_112 | _T_171; // @[Replacement.scala 111:72]
  wire [3:0] _T_175 = _T_173 ? 4'h0 : _T_174; // @[Replacement.scala 111:20]
  wire  _T_176 = 6'h1 == replacerWayWire; // @[Replacement.scala 111:25]
  wire [3:0] _T_177 = _T_114 | _T_171; // @[Replacement.scala 111:72]
  wire [3:0] _T_178 = _T_176 ? 4'h0 : _T_177; // @[Replacement.scala 111:20]
  wire  _T_179 = 6'h2 == replacerWayWire; // @[Replacement.scala 111:25]
  wire [3:0] _T_180 = _T_116 | _T_171; // @[Replacement.scala 111:72]
  wire [3:0] _T_181 = _T_179 ? 4'h0 : _T_180; // @[Replacement.scala 111:20]
  wire [5:0] _T_186 = {_T_181[3],_T_178[3:2],_T_175[3:1]}; // @[Cat.scala 29:58]
  wire  missLD = _T_69; // @[programmableCache.scala 111:22 programmableCache.scala 277:12]
  wire [3:0] tbeWay = input__io_deq_bits_tbeOut_way; // @[programmableCache.scala 294:12]
  wire  _T_187 = tbeWay == 4'h4; // @[programmableCache.scala 363:44]
  reg [3:0] wayInputCache; // @[Reg.scala 27:20]
  reg [31:0] tbeFields_0; // @[Reg.scala 27:20]
  reg [5:0] _T_194; // @[Reg.scala 27:20]
  reg [31:0] inputToPC_addr; // @[Reg.scala 27:20]
  reg [63:0] inputToPC_data; // @[Reg.scala 27:20]
  wire  _T_200 = actionReg_0_io_deq_bits_action_actionType == 4'h0; // @[programmableCache.scala 371:73]
  wire  isCacheAction_0 = _T_200 & actionReg_0_io_deq_valid; // @[programmableCache.scala 371:82]
  wire  _T_202 = actionReg_0_io_deq_bits_action_actionType == 4'h2; // @[programmableCache.scala 372:77]
  wire  _T_206 = actionReg_0_io_deq_bits_action_actionType == 4'h4; // @[programmableCache.scala 374:72]
  wire  _T_208 = actionReg_0_io_deq_bits_action_actionType >= 4'h8; // @[programmableCache.scala 375:73]
  wire [15:0] pcWire_0_pc = pc_io_read_0_out_bits_pc; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [31:0] _GEN_279 = 6'h1 == pcWire_0_pc[5:0] ? 32'h10000001 : 32'h0; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_280 = 6'h2 == pcWire_0_pc[5:0] ? 32'h34 : _GEN_279; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_281 = 6'h3 == pcWire_0_pc[5:0] ? 32'he2000010 : _GEN_280; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_282 = 6'h4 == pcWire_0_pc[5:0] ? 32'h40000203 : _GEN_281; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_283 = 6'h5 == pcWire_0_pc[5:0] ? 32'h20001108 : _GEN_282; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_284 = 6'h6 == pcWire_0_pc[5:0] ? 32'h30000001 : _GEN_283; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_285 = 6'h7 == pcWire_0_pc[5:0] ? 32'h0 : _GEN_284; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_286 = 6'h8 == pcWire_0_pc[5:0] ? 32'hc0000827 : _GEN_285; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_287 = 6'h9 == pcWire_0_pc[5:0] ? 32'h10000000 : _GEN_286; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_288 = 6'ha == pcWire_0_pc[5:0] ? 32'h30000001 : _GEN_287; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_289 = 6'hb == pcWire_0_pc[5:0] ? 32'h0 : _GEN_288; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_290 = 6'hc == pcWire_0_pc[5:0] ? 32'h10000001 : _GEN_289; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_291 = 6'hd == pcWire_0_pc[5:0] ? 32'h34 : _GEN_290; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_292 = 6'he == pcWire_0_pc[5:0] ? 32'h20001108 : _GEN_291; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_293 = 6'hf == pcWire_0_pc[5:0] ? 32'h30000004 : _GEN_292; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_294 = 6'h10 == pcWire_0_pc[5:0] ? 32'h0 : _GEN_293; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_295 = 6'h11 == pcWire_0_pc[5:0] ? 32'h10000002 : _GEN_294; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_296 = 6'h12 == pcWire_0_pc[5:0] ? 32'h80 : _GEN_295; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_297 = 6'h13 == pcWire_0_pc[5:0] ? 32'h100 : _GEN_296; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_298 = 6'h14 == pcWire_0_pc[5:0] ? 32'h30000002 : _GEN_297; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_299 = 6'h15 == pcWire_0_pc[5:0] ? 32'h0 : _GEN_298; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_300 = 6'h16 == pcWire_0_pc[5:0] ? 32'h10000002 : _GEN_299; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_301 = 6'h17 == pcWire_0_pc[5:0] ? 32'h80 : _GEN_300; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_302 = 6'h18 == pcWire_0_pc[5:0] ? 32'h30000002 : _GEN_301; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_303 = 6'h19 == pcWire_0_pc[5:0] ? 32'h0 : _GEN_302; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_304 = 6'h1a == pcWire_0_pc[5:0] ? 32'h20000108 : _GEN_303; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_305 = 6'h1b == pcWire_0_pc[5:0] ? 32'h30000002 : _GEN_304; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_306 = 6'h1c == pcWire_0_pc[5:0] ? 32'h0 : _GEN_305; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_307 = 6'h1d == pcWire_0_pc[5:0] ? 32'h34 : _GEN_306; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_308 = 6'h1e == pcWire_0_pc[5:0] ? 32'h80 : _GEN_307; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_309 = 6'h1f == pcWire_0_pc[5:0] ? 32'h100 : _GEN_308; // @[Gem5CacheLogic.scala 110:53]
  wire [31:0] _GEN_310 = 6'h20 == pcWire_0_pc[5:0] ? 32'h30000002 : _GEN_309; // @[Gem5CacheLogic.scala 110:53]
  wire  _T_223 = pc_io_read_0_out_bits_way == 3'h4; // @[programmableCache.scala 396:52]
  wire  updateWay_0 = _T_223 & cache_io_cpu_0_resp_valid; // @[programmableCache.scala 396:64]
  wire [3:0] cacheWayWire_0 = {{1'd0}, cache_io_cpu_0_resp_bits_way}; // @[programmableCache.scala 154:28 programmableCache.scala 213:25]
  wire [2:0] pcWire_0_way = pc_io_read_0_out_bits_way; // @[programmableCache.scala 116:22 programmableCache.scala 407:19]
  wire [3:0] _T_214 = updateWay_0 ? cacheWayWire_0 : {{1'd0}, pcWire_0_way}; // @[programmableCache.scala 386:45]
  wire  firstLineNextRoutine_0 = _GEN_310 == 32'h0; // @[programmableCache.scala 392:72]
  wire [15:0] _T_218 = pcWire_0_pc + 16'h1; // @[programmableCache.scala 393:81]
  wire [15:0] _T_220 = _T_218 + compUnit_0_io_pc; // @[programmableCache.scala 393:87]
  wire [3:0] _T_225 = updateWay_0 ? cacheWayWire_0 : {{1'd0}, pc_io_read_0_out_bits_way}; // @[programmableCache.scala 398:46]
  wire [31:0] instruction_bits_addr = inputArbiter_io_out_bits_addr; // @[programmableCache.scala 110:27 programmableCache.scala 252:17]
  wire  _T_259 = mimoQ_io_deq_bits_0_way != 3'h4; // @[programmableCache.scala 471:83]
  wire [63:0] _GEN_382 = 2'h1 == actionReg_0_io_deq_bits_action_signals[2:1] ? compUnit_0_io_reg_file_1 : _GEN_377; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_383 = 2'h2 == actionReg_0_io_deq_bits_action_signals[2:1] ? compUnit_0_io_reg_file_2 : _GEN_382; // @[programmableCache.scala 487:47]
  wire [63:0] _GEN_384 = 2'h3 == actionReg_0_io_deq_bits_action_signals[2:1] ? compUnit_0_io_reg_file_3 : _GEN_383; // @[programmableCache.scala 487:47]
  reg [31:0] _T_266; // @[programmableCache.scala 511:55]
  wire  _T_267 = probeWay_io_deq_ready & probeWay_io_deq_valid; // @[Decoupled.scala 40:37]
  reg [1:0] _T_268; // @[programmableCache.scala 531:49]
  reg [31:0] _T_269; // @[programmableCache.scala 531:90]
  reg [63:0] _T_270; // @[programmableCache.scala 531:138]
  wire  _T_272 = ~reset; // @[programmableCache.scala 531:15]
  reg [1:0] _T_273; // @[programmableCache.scala 532:21]
  wire  _T_274 = _T_273 == 2'h3; // @[programmableCache.scala 532:46]
  reg  _T_281; // @[programmableCache.scala 538:31]
  wire  _T_291 = instruction_ready & instruction_valid; // @[Decoupled.scala 40:37]
  wire  _T_294 = _T_52 & _T_74; // @[programmableCache.scala 557:48]
  wire  _T_297 = _T_52 & _T_71; // @[programmableCache.scala 558:48]
  wire  _T_304 = _T_52 & _T_56; // @[programmableCache.scala 559:48]
  wire  hitLD = _T_66; // @[programmableCache.scala 134:29 programmableCache.scala 276:11]
  wire [3:0] replaceWayInputCache = _T_194[3:0]; // @[programmableCache.scala 162:36 programmableCache.scala 365:26]
  wire  _GEN_390 = _T_267 & _T_274; // @[programmableCache.scala 533:19]
  wire  _GEN_392 = _GEN_390 & hitLD; // @[programmableCache.scala 535:23]
  wire  _GEN_394 = ~hitLD; // @[programmableCache.scala 537:23]
  wire  _GEN_395 = _GEN_390 & _GEN_394; // @[programmableCache.scala 537:23]
  wire  _GEN_396 = _GEN_395 & isLocked; // @[programmableCache.scala 537:23]
  wire  _GEN_400 = ~isLocked; // @[programmableCache.scala 539:23]
  wire  _GEN_401 = _GEN_395 & _GEN_400; // @[programmableCache.scala 539:23]
  wire  _GEN_402 = _GEN_401 & _T_281; // @[programmableCache.scala 539:23]
  wire  _GEN_408 = ~_T_281; // @[programmableCache.scala 541:23]
  wire  _GEN_409 = _GEN_401 & _GEN_408; // @[programmableCache.scala 541:23]
  wire  _GEN_410 = _GEN_409 & hit; // @[programmableCache.scala 541:23]
  wire  _GEN_418 = ~hit; // @[programmableCache.scala 543:23]
  wire  _GEN_419 = _GEN_409 & _GEN_418; // @[programmableCache.scala 543:23]
  Gem5Cache cache ( // @[programmableCache.scala 52:26]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_cpu_0_req_valid(cache_io_cpu_0_req_valid),
    .io_cpu_0_req_bits_addr(cache_io_cpu_0_req_bits_addr),
    .io_cpu_0_req_bits_data(cache_io_cpu_0_req_bits_data),
    .io_cpu_0_req_bits_command(cache_io_cpu_0_req_bits_command),
    .io_cpu_0_req_bits_way(cache_io_cpu_0_req_bits_way),
    .io_cpu_0_req_bits_replaceWay(cache_io_cpu_0_req_bits_replaceWay),
    .io_cpu_0_resp_valid(cache_io_cpu_0_resp_valid),
    .io_cpu_0_resp_bits_iswrite(cache_io_cpu_0_resp_bits_iswrite),
    .io_cpu_0_resp_bits_way(cache_io_cpu_0_resp_bits_way),
    .io_probe_req_valid(cache_io_probe_req_valid),
    .io_probe_req_bits_addr(cache_io_probe_req_bits_addr),
    .io_probe_req_bits_command(cache_io_probe_req_bits_command),
    .io_probe_resp_valid(cache_io_probe_resp_valid),
    .io_probe_resp_bits_way(cache_io_probe_resp_bits_way),
    .io_probe_multiWay_valid(cache_io_probe_multiWay_valid),
    .io_probe_multiWay_bits_way_0(cache_io_probe_multiWay_bits_way_0),
    .io_probe_multiWay_bits_way_1(cache_io_probe_multiWay_bits_way_1),
    .io_probe_multiWay_bits_way_2(cache_io_probe_multiWay_bits_way_2),
    .io_probe_multiWay_bits_way_3(cache_io_probe_multiWay_bits_way_3),
    .io_probe_multiWay_bits_addr(cache_io_probe_multiWay_bits_addr),
    .io_bipassLD_in_valid(cache_io_bipassLD_in_valid),
    .io_bipassLD_in_bits_addr(cache_io_bipassLD_in_bits_addr),
    .io_bipassLD_in_bits_way(cache_io_bipassLD_in_bits_way),
    .io_bipassLD_out_valid(cache_io_bipassLD_out_valid),
    .io_bipassLD_out_bits_data(cache_io_bipassLD_out_bits_data)
  );
  TBETable tbe ( // @[programmableCache.scala 53:26]
    .clock(tbe_clock),
    .reset(tbe_reset),
    .io_write_0_valid(tbe_io_write_0_valid),
    .io_write_0_bits_addr(tbe_io_write_0_bits_addr),
    .io_write_0_bits_command(tbe_io_write_0_bits_command),
    .io_write_0_bits_mask(tbe_io_write_0_bits_mask),
    .io_write_0_bits_inputTBE_state_state(tbe_io_write_0_bits_inputTBE_state_state),
    .io_write_0_bits_inputTBE_way(tbe_io_write_0_bits_inputTBE_way),
    .io_write_0_bits_inputTBE_fields_0(tbe_io_write_0_bits_inputTBE_fields_0),
    .io_read_valid(tbe_io_read_valid),
    .io_read_bits_addr(tbe_io_read_bits_addr),
    .io_outputTBE_bits_state_state(tbe_io_outputTBE_bits_state_state),
    .io_outputTBE_bits_way(tbe_io_outputTBE_bits_way),
    .io_outputTBE_bits_fields_0(tbe_io_outputTBE_bits_fields_0),
    .io_isFull(tbe_io_isFull)
  );
  lockVector lockMem ( // @[programmableCache.scala 54:26]
    .clock(lockMem_clock),
    .reset(lockMem_reset),
    .io_lock_in_valid(lockMem_io_lock_in_valid),
    .io_lock_in_bits_addr(lockMem_io_lock_in_bits_addr),
    .io_probe_out_valid(lockMem_io_probe_out_valid),
    .io_probe_out_bits(lockMem_io_probe_out_bits),
    .io_probe_in_valid(lockMem_io_probe_in_valid),
    .io_probe_in_bits_addr(lockMem_io_probe_in_bits_addr),
    .io_unLock_0_in_valid(lockMem_io_unLock_0_in_valid),
    .io_unLock_0_in_bits_addr(lockMem_io_unLock_0_in_bits_addr)
  );
  stateMem stateMem ( // @[programmableCache.scala 55:27]
    .clock(stateMem_clock),
    .reset(stateMem_reset),
    .io_in_0_valid(stateMem_io_in_0_valid),
    .io_in_0_bits_state_state(stateMem_io_in_0_bits_state_state),
    .io_in_0_bits_addr(stateMem_io_in_0_bits_addr),
    .io_in_0_bits_way(stateMem_io_in_0_bits_way),
    .io_in_1_valid(stateMem_io_in_1_valid),
    .io_in_1_bits_addr(stateMem_io_in_1_bits_addr),
    .io_in_1_bits_way(stateMem_io_in_1_bits_way),
    .io_out_valid(stateMem_io_out_valid),
    .io_out_bits_state(stateMem_io_out_bits_state)
  );
  PC pc ( // @[programmableCache.scala 56:26]
    .clock(pc_clock),
    .reset(pc_reset),
    .io_write_ready(pc_io_write_ready),
    .io_write_valid(pc_io_write_valid),
    .io_write_bits_addr(pc_io_write_bits_addr),
    .io_write_bits_way(pc_io_write_bits_way),
    .io_write_bits_data(pc_io_write_bits_data),
    .io_write_bits_replaceWay(pc_io_write_bits_replaceWay),
    .io_write_bits_tbeFields_0(pc_io_write_bits_tbeFields_0),
    .io_write_bits_pc(pc_io_write_bits_pc),
    .io_read_0_in_bits_data_way(pc_io_read_0_in_bits_data_way),
    .io_read_0_in_bits_data_pc(pc_io_read_0_in_bits_data_pc),
    .io_read_0_in_bits_data_valid(pc_io_read_0_in_bits_data_valid),
    .io_read_0_out_bits_addr(pc_io_read_0_out_bits_addr),
    .io_read_0_out_bits_way(pc_io_read_0_out_bits_way),
    .io_read_0_out_bits_data(pc_io_read_0_out_bits_data),
    .io_read_0_out_bits_replaceWay(pc_io_read_0_out_bits_replaceWay),
    .io_read_0_out_bits_tbeFields_0(pc_io_read_0_out_bits_tbeFields_0),
    .io_read_0_out_bits_pc(pc_io_read_0_out_bits_pc),
    .io_read_0_out_bits_valid(pc_io_read_0_out_bits_valid),
    .io_isFull(pc_io_isFull)
  );
  Arbiter_3 inputArbiter ( // @[programmableCache.scala 57:33]
    .io_in_0_valid(inputArbiter_io_in_0_valid),
    .io_in_0_bits_event(inputArbiter_io_in_0_bits_event),
    .io_in_0_bits_addr(inputArbiter_io_in_0_bits_addr),
    .io_in_0_bits_data(inputArbiter_io_in_0_bits_data),
    .io_in_1_ready(inputArbiter_io_in_1_ready),
    .io_in_1_valid(inputArbiter_io_in_1_valid),
    .io_in_1_bits_event(inputArbiter_io_in_1_bits_event),
    .io_in_1_bits_addr(inputArbiter_io_in_1_bits_addr),
    .io_in_1_bits_data(inputArbiter_io_in_1_bits_data),
    .io_in_2_valid(inputArbiter_io_in_2_valid),
    .io_in_2_bits_event(inputArbiter_io_in_2_bits_event),
    .io_in_2_bits_addr(inputArbiter_io_in_2_bits_addr),
    .io_in_2_bits_data(inputArbiter_io_in_2_bits_data),
    .io_in_3_valid(inputArbiter_io_in_3_valid),
    .io_in_3_bits_event(inputArbiter_io_in_3_bits_event),
    .io_in_3_bits_addr(inputArbiter_io_in_3_bits_addr),
    .io_in_3_bits_data(inputArbiter_io_in_3_bits_data),
    .io_out_ready(inputArbiter_io_out_ready),
    .io_out_valid(inputArbiter_io_out_valid),
    .io_out_bits_event(inputArbiter_io_out_bits_event),
    .io_out_bits_addr(inputArbiter_io_out_bits_addr),
    .io_out_bits_data(inputArbiter_io_out_bits_data),
    .io_chosen(inputArbiter_io_chosen)
  );
  RRArbiter_2 outReqArbiter ( // @[programmableCache.scala 58:33]
    .io_in_0_valid(outReqArbiter_io_in_0_valid),
    .io_in_0_bits_req_addr(outReqArbiter_io_in_0_bits_req_addr),
    .io_in_0_bits_req_inst(outReqArbiter_io_in_0_bits_req_inst),
    .io_in_0_bits_req_data(outReqArbiter_io_in_0_bits_req_data),
    .io_out_valid(outReqArbiter_io_out_valid),
    .io_out_bits_req_addr(outReqArbiter_io_out_bits_req_addr),
    .io_out_bits_req_inst(outReqArbiter_io_out_bits_req_inst),
    .io_out_bits_req_data(outReqArbiter_io_out_bits_req_data)
  );
  Arbiter_4 outRespArbiter ( // @[programmableCache.scala 59:33]
    .io_in_0_valid(outRespArbiter_io_in_0_valid),
    .io_in_0_bits_addr(outRespArbiter_io_in_0_bits_addr),
    .io_in_1_valid(outRespArbiter_io_in_1_valid),
    .io_in_1_bits_addr(outRespArbiter_io_in_1_bits_addr),
    .io_out_valid(outRespArbiter_io_out_valid),
    .io_out_bits_addr(outRespArbiter_io_out_bits_addr)
  );
  Arbiter_5 feedbackArbiter ( // @[programmableCache.scala 60:34]
    .io_in_0_ready(feedbackArbiter_io_in_0_ready),
    .io_in_0_valid(feedbackArbiter_io_in_0_valid),
    .io_in_0_bits_event(feedbackArbiter_io_in_0_bits_event),
    .io_in_0_bits_addr(feedbackArbiter_io_in_0_bits_addr),
    .io_in_0_bits_data(feedbackArbiter_io_in_0_bits_data),
    .io_out_ready(feedbackArbiter_io_out_ready),
    .io_out_valid(feedbackArbiter_io_out_valid),
    .io_out_bits_event(feedbackArbiter_io_out_bits_event),
    .io_out_bits_addr(feedbackArbiter_io_out_bits_addr),
    .io_out_bits_data(feedbackArbiter_io_out_bits_data)
  );
  Queue_7 input_ ( // @[programmableCache.scala 90:23]
    .clock(input__clock),
    .reset(input__reset),
    .io_enq_ready(input__io_enq_ready),
    .io_enq_valid(input__io_enq_valid),
    .io_enq_bits_inst_event(input__io_enq_bits_inst_event),
    .io_enq_bits_inst_addr(input__io_enq_bits_inst_addr),
    .io_enq_bits_inst_data(input__io_enq_bits_inst_data),
    .io_enq_bits_tbeOut_state_state(input__io_enq_bits_tbeOut_state_state),
    .io_enq_bits_tbeOut_way(input__io_enq_bits_tbeOut_way),
    .io_enq_bits_tbeOut_fields_0(input__io_enq_bits_tbeOut_fields_0),
    .io_deq_ready(input__io_deq_ready),
    .io_deq_valid(input__io_deq_valid),
    .io_deq_bits_inst_event(input__io_deq_bits_inst_event),
    .io_deq_bits_inst_addr(input__io_deq_bits_inst_addr),
    .io_deq_bits_inst_data(input__io_deq_bits_inst_data),
    .io_deq_bits_tbeOut_state_state(input__io_deq_bits_tbeOut_state_state),
    .io_deq_bits_tbeOut_way(input__io_deq_bits_tbeOut_way),
    .io_deq_bits_tbeOut_fields_0(input__io_deq_bits_tbeOut_fields_0)
  );
  Queue_8 respPortQueue_0 ( // @[programmableCache.scala 93:27]
    .clock(respPortQueue_0_clock),
    .reset(respPortQueue_0_reset),
    .io_enq_ready(respPortQueue_0_io_enq_ready),
    .io_enq_valid(respPortQueue_0_io_enq_valid),
    .io_enq_bits_event(respPortQueue_0_io_enq_bits_event),
    .io_enq_bits_addr(respPortQueue_0_io_enq_bits_addr),
    .io_enq_bits_data(respPortQueue_0_io_enq_bits_data),
    .io_deq_ready(respPortQueue_0_io_deq_ready),
    .io_deq_valid(respPortQueue_0_io_deq_valid),
    .io_deq_bits_event(respPortQueue_0_io_deq_bits_event),
    .io_deq_bits_addr(respPortQueue_0_io_deq_bits_addr),
    .io_deq_bits_data(respPortQueue_0_io_deq_bits_data)
  );
  Queue_8 respPortQueue_1 ( // @[programmableCache.scala 93:27]
    .clock(respPortQueue_1_clock),
    .reset(respPortQueue_1_reset),
    .io_enq_ready(respPortQueue_1_io_enq_ready),
    .io_enq_valid(respPortQueue_1_io_enq_valid),
    .io_enq_bits_event(respPortQueue_1_io_enq_bits_event),
    .io_enq_bits_addr(respPortQueue_1_io_enq_bits_addr),
    .io_enq_bits_data(respPortQueue_1_io_enq_bits_data),
    .io_deq_ready(respPortQueue_1_io_deq_ready),
    .io_deq_valid(respPortQueue_1_io_deq_valid),
    .io_deq_bits_event(respPortQueue_1_io_deq_bits_event),
    .io_deq_bits_addr(respPortQueue_1_io_deq_bits_addr),
    .io_deq_bits_data(respPortQueue_1_io_deq_bits_data)
  );
  Queue_10 reqPortQueue_0 ( // @[programmableCache.scala 98:27]
    .clock(reqPortQueue_0_clock),
    .reset(reqPortQueue_0_reset),
    .io_enq_ready(reqPortQueue_0_io_enq_ready),
    .io_enq_valid(reqPortQueue_0_io_enq_valid),
    .io_enq_bits_addr(reqPortQueue_0_io_enq_bits_addr),
    .io_enq_bits_data(reqPortQueue_0_io_enq_bits_data),
    .io_deq_valid(reqPortQueue_0_io_deq_valid),
    .io_deq_bits_addr(reqPortQueue_0_io_deq_bits_addr),
    .io_deq_bits_inst(reqPortQueue_0_io_deq_bits_inst),
    .io_deq_bits_data(reqPortQueue_0_io_deq_bits_data)
  );
  Queue_8 feedbackInQueue_0 ( // @[programmableCache.scala 104:27]
    .clock(feedbackInQueue_0_clock),
    .reset(feedbackInQueue_0_reset),
    .io_enq_ready(feedbackInQueue_0_io_enq_ready),
    .io_enq_valid(feedbackInQueue_0_io_enq_valid),
    .io_enq_bits_event(feedbackInQueue_0_io_enq_bits_event),
    .io_enq_bits_addr(feedbackInQueue_0_io_enq_bits_addr),
    .io_enq_bits_data(feedbackInQueue_0_io_enq_bits_data),
    .io_deq_ready(feedbackInQueue_0_io_deq_ready),
    .io_deq_valid(feedbackInQueue_0_io_deq_valid),
    .io_deq_bits_event(feedbackInQueue_0_io_deq_bits_event),
    .io_deq_bits_addr(feedbackInQueue_0_io_deq_bits_addr),
    .io_deq_bits_data(feedbackInQueue_0_io_deq_bits_data)
  );
  Queue_12 probeWay ( // @[programmableCache.scala 108:26]
    .clock(probeWay_clock),
    .reset(probeWay_reset),
    .io_enq_ready(probeWay_io_enq_ready),
    .io_enq_valid(probeWay_io_enq_valid),
    .io_enq_bits(probeWay_io_enq_bits),
    .io_deq_ready(probeWay_io_deq_ready),
    .io_deq_valid(probeWay_io_deq_valid),
    .io_deq_bits(probeWay_io_deq_bits)
  );
  Queue_8 feedbackOutQueue ( // @[programmableCache.scala 165:34]
    .clock(feedbackOutQueue_clock),
    .reset(feedbackOutQueue_reset),
    .io_enq_ready(feedbackOutQueue_io_enq_ready),
    .io_enq_valid(feedbackOutQueue_io_enq_valid),
    .io_enq_bits_event(feedbackOutQueue_io_enq_bits_event),
    .io_enq_bits_addr(feedbackOutQueue_io_enq_bits_addr),
    .io_enq_bits_data(feedbackOutQueue_io_enq_bits_data),
    .io_deq_ready(feedbackOutQueue_io_deq_ready),
    .io_deq_valid(feedbackOutQueue_io_deq_valid),
    .io_deq_bits_event(feedbackOutQueue_io_deq_bits_event),
    .io_deq_bits_addr(feedbackOutQueue_io_deq_bits_addr),
    .io_deq_bits_data(feedbackOutQueue_io_deq_bits_data)
  );
  Queue_14 routineQueue ( // @[programmableCache.scala 166:30]
    .clock(routineQueue_clock),
    .reset(routineQueue_reset),
    .io_enq_ready(routineQueue_io_enq_ready),
    .io_enq_valid(routineQueue_io_enq_valid),
    .io_enq_bits(routineQueue_io_enq_bits),
    .io_deq_ready(routineQueue_io_deq_ready),
    .io_deq_valid(routineQueue_io_deq_valid),
    .io_deq_bits(routineQueue_io_deq_bits)
  );
  Queue_15 actionReg_0 ( // @[programmableCache.scala 169:32]
    .clock(actionReg_0_clock),
    .reset(actionReg_0_reset),
    .io_enq_ready(actionReg_0_io_enq_ready),
    .io_enq_valid(actionReg_0_io_enq_valid),
    .io_enq_bits_addr(actionReg_0_io_enq_bits_addr),
    .io_enq_bits_way(actionReg_0_io_enq_bits_way),
    .io_enq_bits_data(actionReg_0_io_enq_bits_data),
    .io_enq_bits_replaceWay(actionReg_0_io_enq_bits_replaceWay),
    .io_enq_bits_tbeFields_0(actionReg_0_io_enq_bits_tbeFields_0),
    .io_enq_bits_action_signals(actionReg_0_io_enq_bits_action_signals),
    .io_enq_bits_action_actionType(actionReg_0_io_enq_bits_action_actionType),
    .io_deq_ready(actionReg_0_io_deq_ready),
    .io_deq_valid(actionReg_0_io_deq_valid),
    .io_deq_bits_addr(actionReg_0_io_deq_bits_addr),
    .io_deq_bits_way(actionReg_0_io_deq_bits_way),
    .io_deq_bits_data(actionReg_0_io_deq_bits_data),
    .io_deq_bits_replaceWay(actionReg_0_io_deq_bits_replaceWay),
    .io_deq_bits_tbeFields_0(actionReg_0_io_deq_bits_tbeFields_0),
    .io_deq_bits_action_signals(actionReg_0_io_deq_bits_action_signals),
    .io_deq_bits_action_actionType(actionReg_0_io_deq_bits_action_actionType)
  );
  MIMOQueue mimoQ ( // @[programmableCache.scala 173:24]
    .clock(mimoQ_clock),
    .reset(mimoQ_reset),
    .io_enq_ready(mimoQ_io_enq_ready),
    .io_enq_valid(mimoQ_io_enq_valid),
    .io_enq_bits_0_way(mimoQ_io_enq_bits_0_way),
    .io_enq_bits_0_addr(mimoQ_io_enq_bits_0_addr),
    .io_enq_bits_1_way(mimoQ_io_enq_bits_1_way),
    .io_enq_bits_1_addr(mimoQ_io_enq_bits_1_addr),
    .io_enq_bits_2_way(mimoQ_io_enq_bits_2_way),
    .io_enq_bits_2_addr(mimoQ_io_enq_bits_2_addr),
    .io_enq_bits_3_way(mimoQ_io_enq_bits_3_way),
    .io_enq_bits_3_addr(mimoQ_io_enq_bits_3_addr),
    .io_deq_valid(mimoQ_io_deq_valid),
    .io_deq_bits_0_way(mimoQ_io_deq_bits_0_way),
    .io_deq_bits_0_addr(mimoQ_io_deq_bits_0_addr),
    .io_count(mimoQ_io_count)
  );
  Computation compUnit_0 ( // @[programmableCache.scala 177:27]
    .clock(compUnit_0_clock),
    .reset(compUnit_0_reset),
    .io_instruction_valid(compUnit_0_io_instruction_valid),
    .io_instruction_bits(compUnit_0_io_instruction_bits),
    .io_clear(compUnit_0_io_clear),
    .io_op1_valid(compUnit_0_io_op1_valid),
    .io_op1_bits(compUnit_0_io_op1_bits),
    .io_op2_valid(compUnit_0_io_op2_valid),
    .io_op2_bits(compUnit_0_io_op2_bits),
    .io_pc(compUnit_0_io_pc),
    .io_reg_file_0(compUnit_0_io_reg_file_0),
    .io_reg_file_1(compUnit_0_io_reg_file_1),
    .io_reg_file_2(compUnit_0_io_reg_file_2),
    .io_reg_file_3(compUnit_0_io_reg_file_3)
  );
  Mux3 compUnitInput1_0 ( // @[programmableCache.scala 182:30]
    .io_in_hardCoded(compUnitInput1_0_io_in_hardCoded),
    .io_in_data(compUnitInput1_0_io_in_data),
    .io_in_tbe(compUnitInput1_0_io_in_tbe),
    .io_in_select(compUnitInput1_0_io_in_select),
    .io_out_valid(compUnitInput1_0_io_out_valid),
    .io_out_bits(compUnitInput1_0_io_out_bits)
  );
  Mux3 compUnitInput2_0 ( // @[programmableCache.scala 188:30]
    .io_in_hardCoded(compUnitInput2_0_io_in_hardCoded),
    .io_in_data(compUnitInput2_0_io_in_data),
    .io_in_tbe(compUnitInput2_0_io_in_tbe),
    .io_in_select(compUnitInput2_0_io_in_select),
    .io_out_valid(compUnitInput2_0_io_out_valid),
    .io_out_bits(compUnitInput2_0_io_out_bits)
  );
  assign io_in_cpu_ready = _T_52 & _T_74; // @[programmableCache.scala 240:37 programmableCache.scala 280:28]
  assign io_in_memCtrl_ready = _T_52 & _T_71; // @[programmableCache.scala 241:41 programmableCache.scala 279:28]
  assign io_in_otherNodes_ready = _T_52 & _T_77; // @[programmableCache.scala 239:44 programmableCache.scala 281:28]
  assign io_out_req_valid = outReqArbiter_io_out_valid; // @[programmableCache.scala 499:22]
  assign io_out_req_bits_req_addr = outReqArbiter_io_out_bits_req_addr; // @[programmableCache.scala 497:30]
  assign io_out_req_bits_req_inst = outReqArbiter_io_out_bits_req_inst; // @[programmableCache.scala 495:30]
  assign io_out_req_bits_req_data = outReqArbiter_io_out_bits_req_data; // @[programmableCache.scala 496:30]
  assign io_out_resp_valid = outRespArbiter_io_out_valid; // @[programmableCache.scala 525:27]
  assign io_out_resp_bits_addr = outRespArbiter_io_out_bits_addr; // @[programmableCache.scala 524:27]
  assign _T_297_0 = _T_72;
  assign _T_291_0 = _T_52;
  assign _T_304_0 = probeStart;
  assign hitLD_0 = hitLD;
  assign missLD_0 = missLD;
  assign _T_294_0 = _T_75;
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_cpu_0_req_valid = actionReg_0_io_deq_ready & actionReg_0_io_deq_valid; // @[programmableCache.scala 460:35]
  assign cache_io_cpu_0_req_bits_addr = actionReg_0_io_deq_bits_addr; // @[programmableCache.scala 459:39]
  assign cache_io_cpu_0_req_bits_data = actionReg_0_io_deq_bits_data; // @[programmableCache.scala 461:39]
  assign cache_io_cpu_0_req_bits_command = isCacheAction_0 ? actionReg_0_io_deq_bits_action_signals : 28'h0; // @[programmableCache.scala 458:42]
  assign cache_io_cpu_0_req_bits_way = actionReg_0_io_deq_bits_way; // @[programmableCache.scala 457:38]
  assign cache_io_cpu_0_req_bits_replaceWay = actionReg_0_io_deq_bits_replaceWay; // @[programmableCache.scala 462:45]
  assign cache_io_probe_req_valid = _T_52 & _T_56; // @[programmableCache.scala 468:30]
  assign cache_io_probe_req_bits_addr = probeStart ? instruction_bits_addr : 32'h0; // @[programmableCache.scala 466:34]
  assign cache_io_probe_req_bits_command = probeStart ? 28'hb : 28'h0; // @[programmableCache.scala 465:37]
  assign cache_io_bipassLD_in_valid = mimoQ_io_deq_valid & _T_259; // @[programmableCache.scala 471:32]
  assign cache_io_bipassLD_in_bits_addr = mimoQ_io_deq_bits_0_addr; // @[programmableCache.scala 472:37]
  assign cache_io_bipassLD_in_bits_way = {{1'd0}, mimoQ_io_deq_bits_0_way}; // @[programmableCache.scala 473:35]
  assign tbe_clock = clock;
  assign tbe_reset = reset;
  assign tbe_io_write_0_valid = isTBEAction_0 | isStateAction_0; // @[programmableCache.scala 309:31]
  assign tbe_io_write_0_bits_addr = {{32'd0}, actionReg_0_io_deq_bits_addr}; // @[programmableCache.scala 306:35]
  assign tbe_io_write_0_bits_command = isStateAction_0 ? 2'h3 : tbeAction_0; // @[programmableCache.scala 305:38]
  assign tbe_io_write_0_bits_mask = isStateAction_0 | maskField_0; // @[programmableCache.scala 308:35]
  assign tbe_io_write_0_bits_inputTBE_state_state = isStateAction_0 ? tbeAction_0 : 2'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_write_0_bits_inputTBE_way = {{1'd0}, actionReg_0_io_deq_bits_way}; // @[programmableCache.scala 307:39]
  assign tbe_io_write_0_bits_inputTBE_fields_0 = _T_98 ? tbeFieldUpdateSrc_0 : 32'h0; // @[programmableCache.scala 307:39]
  assign tbe_io_read_valid = inputArbiter_io_out_valid; // @[programmableCache.scala 297:23]
  assign tbe_io_read_bits_addr = {{32'd0}, inputArbiter_io_out_bits_addr}; // @[programmableCache.scala 298:27]
  assign lockMem_clock = clock;
  assign lockMem_reset = reset;
  assign lockMem_io_lock_in_valid = instruction_ready & instruction_valid; // @[programmableCache.scala 320:35]
  assign lockMem_io_lock_in_bits_addr = inputArbiter_io_out_bits_addr; // @[programmableCache.scala 319:35]
  assign lockMem_io_probe_in_valid = inputArbiter_io_out_valid; // @[programmableCache.scala 315:35]
  assign lockMem_io_probe_in_bits_addr = inputArbiter_io_out_bits_addr; // @[programmableCache.scala 314:35]
  assign lockMem_io_unLock_0_in_valid = _T_204 & actionReg_0_io_deq_valid; // @[programmableCache.scala 328:39]
  assign lockMem_io_unLock_0_in_bits_addr = actionReg_0_io_deq_bits_addr; // @[programmableCache.scala 326:43]
  assign stateMem_clock = clock;
  assign stateMem_reset = reset;
  assign stateMem_io_in_0_valid = _T_204 & actionReg_0_io_deq_valid; // @[programmableCache.scala 338:33]
  assign stateMem_io_in_0_bits_state_state = isStateAction_0 ? tbeAction_0 : 2'h0; // @[programmableCache.scala 336:38]
  assign stateMem_io_in_0_bits_addr = actionReg_0_io_deq_bits_addr; // @[programmableCache.scala 335:37]
  assign stateMem_io_in_0_bits_way = actionReg_0_io_deq_bits_way; // @[programmableCache.scala 337:36]
  assign stateMem_io_in_1_valid = input__io_deq_ready & input__io_deq_valid; // @[programmableCache.scala 345:34]
  assign stateMem_io_in_1_bits_addr = input__io_deq_bits_inst_addr; // @[programmableCache.scala 342:38]
  assign stateMem_io_in_1_bits_way = probeWay_io_deq_bits; // @[programmableCache.scala 344:37]
  assign pc_clock = clock;
  assign pc_reset = reset;
  assign pc_io_write_valid = routineQueue_io_deq_ready & routineQueue_io_deq_valid; // @[programmableCache.scala 451:23]
  assign pc_io_write_bits_addr = inputToPC_addr; // @[programmableCache.scala 443:27]
  assign pc_io_write_bits_way = wayInputCache[2:0]; // @[programmableCache.scala 444:26]
  assign pc_io_write_bits_data = inputToPC_data; // @[programmableCache.scala 448:27]
  assign pc_io_write_bits_replaceWay = replaceWayInputCache[2:0]; // @[programmableCache.scala 446:33]
  assign pc_io_write_bits_tbeFields_0 = tbeFields_0; // @[programmableCache.scala 445:32]
  assign pc_io_write_bits_pc = routineQueue_io_deq_bits; // @[programmableCache.scala 447:25]
  assign pc_io_read_0_in_bits_data_way = _T_225[2:0]; // @[programmableCache.scala 398:40]
  assign pc_io_read_0_in_bits_data_pc = firstLineNextRoutine_0 ? pcWire_0_pc : _T_220; // @[programmableCache.scala 400:39]
  assign pc_io_read_0_in_bits_data_valid = ~firstLineNextRoutine_0; // @[programmableCache.scala 403:42]
  assign inputArbiter_io_in_0_valid = io_in_memCtrl_valid; // @[programmableCache.scala 241:41]
  assign inputArbiter_io_in_0_bits_event = io_in_memCtrl_bits_event; // @[programmableCache.scala 241:41]
  assign inputArbiter_io_in_0_bits_addr = io_in_memCtrl_bits_addr; // @[programmableCache.scala 241:41]
  assign inputArbiter_io_in_0_bits_data = io_in_memCtrl_bits_data; // @[programmableCache.scala 241:41]
  assign inputArbiter_io_in_1_valid = feedbackOutQueue_io_deq_valid; // @[programmableCache.scala 242:42]
  assign inputArbiter_io_in_1_bits_event = feedbackOutQueue_io_deq_bits_event; // @[programmableCache.scala 242:42]
  assign inputArbiter_io_in_1_bits_addr = feedbackOutQueue_io_deq_bits_addr; // @[programmableCache.scala 242:42]
  assign inputArbiter_io_in_1_bits_data = feedbackOutQueue_io_deq_bits_data; // @[programmableCache.scala 242:42]
  assign inputArbiter_io_in_2_valid = io_in_otherNodes_valid; // @[programmableCache.scala 239:44]
  assign inputArbiter_io_in_2_bits_event = io_in_otherNodes_bits_event; // @[programmableCache.scala 239:44]
  assign inputArbiter_io_in_2_bits_addr = io_in_otherNodes_bits_addr; // @[programmableCache.scala 239:44]
  assign inputArbiter_io_in_2_bits_data = io_in_otherNodes_bits_data; // @[programmableCache.scala 239:44]
  assign inputArbiter_io_in_3_valid = io_in_cpu_valid; // @[programmableCache.scala 240:37]
  assign inputArbiter_io_in_3_bits_event = io_in_cpu_bits_event; // @[programmableCache.scala 240:37]
  assign inputArbiter_io_in_3_bits_addr = io_in_cpu_bits_addr; // @[programmableCache.scala 240:37]
  assign inputArbiter_io_in_3_bits_data = io_in_cpu_bits_data; // @[programmableCache.scala 240:37]
  assign inputArbiter_io_out_ready = _T_85 & _T_86; // @[programmableCache.scala 252:17]
  assign outReqArbiter_io_in_0_valid = reqPortQueue_0_io_deq_valid; // @[programmableCache.scala 481:41]
  assign outReqArbiter_io_in_0_bits_req_addr = reqPortQueue_0_io_deq_bits_addr; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_0_bits_req_inst = reqPortQueue_0_io_deq_bits_inst; // @[programmableCache.scala 479:41]
  assign outReqArbiter_io_in_0_bits_req_data = reqPortQueue_0_io_deq_bits_data; // @[programmableCache.scala 479:41]
  assign outRespArbiter_io_in_0_valid = respPortQueue_0_io_deq_valid; // @[programmableCache.scala 518:44]
  assign outRespArbiter_io_in_0_bits_addr = respPortQueue_0_io_deq_bits_addr; // @[programmableCache.scala 517:44]
  assign outRespArbiter_io_in_1_valid = respPortQueue_1_io_deq_valid; // @[programmableCache.scala 518:44]
  assign outRespArbiter_io_in_1_bits_addr = respPortQueue_1_io_deq_bits_addr; // @[programmableCache.scala 517:44]
  assign feedbackArbiter_io_in_0_valid = feedbackInQueue_0_io_deq_valid; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_0_bits_event = feedbackInQueue_0_io_deq_bits_event; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_0_bits_addr = feedbackInQueue_0_io_deq_bits_addr; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_in_0_bits_data = feedbackInQueue_0_io_deq_bits_data; // @[programmableCache.scala 246:34]
  assign feedbackArbiter_io_out_ready = feedbackOutQueue_io_enq_ready; // @[programmableCache.scala 244:29]
  assign input__clock = clock;
  assign input__reset = reset;
  assign input__io_enq_valid = _T_91 & _T_86; // @[programmableCache.scala 286:24]
  assign input__io_enq_bits_inst_event = inputArbiter_io_out_bits_event; // @[programmableCache.scala 288:28]
  assign input__io_enq_bits_inst_addr = inputArbiter_io_out_bits_addr; // @[programmableCache.scala 288:28]
  assign input__io_enq_bits_inst_data = inputArbiter_io_out_bits_data; // @[programmableCache.scala 288:28]
  assign input__io_enq_bits_tbeOut_state_state = tbe_io_outputTBE_bits_state_state; // @[programmableCache.scala 289:30]
  assign input__io_enq_bits_tbeOut_way = tbe_io_outputTBE_bits_way; // @[programmableCache.scala 289:30]
  assign input__io_enq_bits_tbeOut_fields_0 = tbe_io_outputTBE_bits_fields_0; // @[programmableCache.scala 289:30]
  assign input__io_deq_ready = routineQueue_io_enq_ready; // @[programmableCache.scala 351:24]
  assign respPortQueue_0_clock = clock;
  assign respPortQueue_0_reset = reset;
  assign respPortQueue_0_io_enq_valid = cache_io_cpu_0_resp_valid & cache_io_cpu_0_resp_bits_iswrite; // @[programmableCache.scala 506:44]
  assign respPortQueue_0_io_enq_bits_event = 2'h0; // @[programmableCache.scala 504:44]
  assign respPortQueue_0_io_enq_bits_addr = actionReg_0_io_deq_bits_addr; // @[programmableCache.scala 505:44]
  assign respPortQueue_0_io_enq_bits_data = 64'h0; // @[programmableCache.scala 503:44]
  assign respPortQueue_0_io_deq_ready = 1'h1; // @[programmableCache.scala 519:39]
  assign respPortQueue_1_clock = clock;
  assign respPortQueue_1_reset = reset;
  assign respPortQueue_1_io_enq_valid = cache_io_bipassLD_out_valid; // @[programmableCache.scala 512:45]
  assign respPortQueue_1_io_enq_bits_event = 2'h0; // @[programmableCache.scala 510:45]
  assign respPortQueue_1_io_enq_bits_addr = _T_266; // @[programmableCache.scala 511:45]
  assign respPortQueue_1_io_enq_bits_data = cache_io_bipassLD_out_bits_data; // @[programmableCache.scala 509:45]
  assign respPortQueue_1_io_deq_ready = 1'h1; // @[programmableCache.scala 519:39]
  assign reqPortQueue_0_clock = clock;
  assign reqPortQueue_0_reset = reset;
  assign reqPortQueue_0_io_enq_valid = _T_206 & actionReg_0_io_deq_valid; // @[programmableCache.scala 490:38]
  assign reqPortQueue_0_io_enq_bits_addr = actionReg_0_io_deq_bits_addr; // @[programmableCache.scala 488:42]
  assign reqPortQueue_0_io_enq_bits_data = actionReg_0_io_deq_bits_action_signals[0] ? _GEN_384 : {{32'd0}, actionReg_0_io_deq_bits_addr}; // @[programmableCache.scala 487:41]
  assign feedbackInQueue_0_clock = clock;
  assign feedbackInQueue_0_reset = reset;
  assign feedbackInQueue_0_io_enq_valid = _T_202 & actionReg_0_io_deq_valid; // @[programmableCache.scala 250:41]
  assign feedbackInQueue_0_io_enq_bits_event = actionReg_0_io_deq_bits_action_signals[13:12]; // @[programmableCache.scala 248:46]
  assign feedbackInQueue_0_io_enq_bits_addr = actionReg_0_io_deq_bits_addr + _GEN_385; // @[programmableCache.scala 247:45]
  assign feedbackInQueue_0_io_enq_bits_data = actionReg_0_io_deq_bits_data - _GEN_386; // @[programmableCache.scala 249:45]
  assign feedbackInQueue_0_io_deq_ready = feedbackArbiter_io_in_0_ready; // @[programmableCache.scala 246:34]
  assign probeWay_clock = clock;
  assign probeWay_reset = reset;
  assign probeWay_io_enq_valid = cache_io_probe_resp_valid; // @[programmableCache.scala 217:29]
  assign probeWay_io_enq_bits = cache_io_probe_resp_bits_way; // @[programmableCache.scala 216:28]
  assign probeWay_io_deq_ready = input__io_deq_ready & input__io_deq_valid; // @[programmableCache.scala 227:29]
  assign feedbackOutQueue_clock = clock;
  assign feedbackOutQueue_reset = reset;
  assign feedbackOutQueue_io_enq_valid = feedbackArbiter_io_out_valid; // @[programmableCache.scala 244:29]
  assign feedbackOutQueue_io_enq_bits_event = feedbackArbiter_io_out_bits_event; // @[programmableCache.scala 244:29]
  assign feedbackOutQueue_io_enq_bits_addr = feedbackArbiter_io_out_bits_addr; // @[programmableCache.scala 244:29]
  assign feedbackOutQueue_io_enq_bits_data = feedbackArbiter_io_out_bits_data; // @[programmableCache.scala 244:29]
  assign feedbackOutQueue_io_deq_ready = inputArbiter_io_in_1_ready; // @[programmableCache.scala 242:42]
  assign routineQueue_clock = clock;
  assign routineQueue_reset = reset;
  assign routineQueue_io_enq_valid = input__io_deq_valid; // @[programmableCache.scala 350:31]
  assign routineQueue_io_enq_bits = {{11'd0}, _GEN_15}; // @[programmableCache.scala 349:30]
  assign routineQueue_io_deq_ready = ~pc_io_isFull; // @[programmableCache.scala 352:31]
  assign actionReg_0_clock = clock;
  assign actionReg_0_reset = reset;
  assign actionReg_0_io_enq_valid = pc_io_read_0_out_bits_valid; // @[programmableCache.scala 438:35]
  assign actionReg_0_io_enq_bits_addr = pc_io_read_0_out_bits_addr; // @[programmableCache.scala 385:39]
  assign actionReg_0_io_enq_bits_way = _T_214[2:0]; // @[programmableCache.scala 386:39]
  assign actionReg_0_io_enq_bits_data = pc_io_read_0_out_bits_data; // @[programmableCache.scala 387:39]
  assign actionReg_0_io_enq_bits_replaceWay = pc_io_read_0_out_bits_replaceWay; // @[programmableCache.scala 388:45]
  assign actionReg_0_io_enq_bits_tbeFields_0 = pc_io_read_0_out_bits_tbeFields_0; // @[programmableCache.scala 390:44]
  assign actionReg_0_io_enq_bits_action_signals = _GEN_310[27:0]; // @[programmableCache.scala 383:49]
  assign actionReg_0_io_enq_bits_action_actionType = _GEN_310[31:28]; // @[programmableCache.scala 384:52]
  assign actionReg_0_io_deq_ready = 1'h1; // @[programmableCache.scala 437:35]
  assign mimoQ_clock = clock;
  assign mimoQ_reset = reset;
  assign mimoQ_io_enq_valid = cache_io_probe_multiWay_valid; // @[programmableCache.scala 222:24]
  assign mimoQ_io_enq_bits_0_way = cache_io_probe_multiWay_bits_way_0; // @[programmableCache.scala 219:56]
  assign mimoQ_io_enq_bits_0_addr = cache_io_probe_multiWay_bits_addr; // @[programmableCache.scala 220:57]
  assign mimoQ_io_enq_bits_1_way = cache_io_probe_multiWay_bits_way_1; // @[programmableCache.scala 219:56]
  assign mimoQ_io_enq_bits_1_addr = cache_io_probe_multiWay_bits_addr; // @[programmableCache.scala 220:57]
  assign mimoQ_io_enq_bits_2_way = cache_io_probe_multiWay_bits_way_2; // @[programmableCache.scala 219:56]
  assign mimoQ_io_enq_bits_2_addr = cache_io_probe_multiWay_bits_addr; // @[programmableCache.scala 220:57]
  assign mimoQ_io_enq_bits_3_way = cache_io_probe_multiWay_bits_way_3; // @[programmableCache.scala 219:56]
  assign mimoQ_io_enq_bits_3_addr = cache_io_probe_multiWay_bits_addr; // @[programmableCache.scala 220:57]
  assign compUnit_0_clock = clock;
  assign compUnit_0_reset = reset;
  assign compUnit_0_io_instruction_valid = _T_208 & actionReg_0_io_deq_valid; // @[programmableCache.scala 435:42]
  assign compUnit_0_io_instruction_bits = actionReg_0_io_deq_bits_action_signals; // @[programmableCache.scala 434:41]
  assign compUnit_0_io_clear = _T_204 & actionReg_0_io_deq_valid; // @[programmableCache.scala 381:30]
  assign compUnit_0_io_op1_valid = compUnitInput1_0_io_out_valid; // @[programmableCache.scala 425:28]
  assign compUnit_0_io_op1_bits = compUnitInput1_0_io_out_bits; // @[programmableCache.scala 425:28]
  assign compUnit_0_io_op2_valid = compUnitInput2_0_io_out_valid; // @[programmableCache.scala 432:28]
  assign compUnit_0_io_op2_bits = compUnitInput2_0_io_out_bits; // @[programmableCache.scala 432:28]
  assign compUnitInput1_0_io_in_hardCoded = 64'h0;
  assign compUnitInput1_0_io_in_data = 64'h0;
  assign compUnitInput1_0_io_in_tbe = {{32'd0}, actionReg_0_io_deq_bits_addr}; // @[programmableCache.scala 422:38]
  assign compUnitInput1_0_io_in_select = {{1'd0}, actionReg_0_io_deq_bits_action_actionType[0]}; // @[programmableCache.scala 424:40]
  assign compUnitInput2_0_io_in_hardCoded = {{48'd0}, actionReg_0_io_deq_bits_action_signals[27:12]}; // @[programmableCache.scala 430:43]
  assign compUnitInput2_0_io_in_data = actionReg_0_io_deq_bits_data; // @[programmableCache.scala 428:38]
  assign compUnitInput2_0_io_in_tbe = {{32'd0}, actionReg_0_io_deq_bits_tbeFields_0}; // @[programmableCache.scala 429:38]
  assign compUnitInput2_0_io_in_select = actionReg_0_io_deq_bits_action_actionType[2:1]; // @[programmableCache.scala 431:40]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  instUsed = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  replStateReg_0 = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  replStateReg_1 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  replStateReg_2 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  replStateReg_3 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  replStateReg_4 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  replStateReg_5 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  replStateReg_6 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  replStateReg_7 = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  replStateReg_8 = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  replStateReg_9 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  replStateReg_10 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  replStateReg_11 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  replStateReg_12 = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  replStateReg_13 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  replStateReg_14 = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  replStateReg_15 = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  replStateReg_16 = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  replStateReg_17 = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  replStateReg_18 = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  replStateReg_19 = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  replStateReg_20 = _RAND_21[5:0];
  _RAND_22 = {1{`RANDOM}};
  replStateReg_21 = _RAND_22[5:0];
  _RAND_23 = {1{`RANDOM}};
  replStateReg_22 = _RAND_23[5:0];
  _RAND_24 = {1{`RANDOM}};
  replStateReg_23 = _RAND_24[5:0];
  _RAND_25 = {1{`RANDOM}};
  replStateReg_24 = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  replStateReg_25 = _RAND_26[5:0];
  _RAND_27 = {1{`RANDOM}};
  replStateReg_26 = _RAND_27[5:0];
  _RAND_28 = {1{`RANDOM}};
  replStateReg_27 = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  replStateReg_28 = _RAND_29[5:0];
  _RAND_30 = {1{`RANDOM}};
  replStateReg_29 = _RAND_30[5:0];
  _RAND_31 = {1{`RANDOM}};
  replStateReg_30 = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  replStateReg_31 = _RAND_32[5:0];
  _RAND_33 = {1{`RANDOM}};
  replStateReg_32 = _RAND_33[5:0];
  _RAND_34 = {1{`RANDOM}};
  replStateReg_33 = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  replStateReg_34 = _RAND_35[5:0];
  _RAND_36 = {1{`RANDOM}};
  replStateReg_35 = _RAND_36[5:0];
  _RAND_37 = {1{`RANDOM}};
  replStateReg_36 = _RAND_37[5:0];
  _RAND_38 = {1{`RANDOM}};
  replStateReg_37 = _RAND_38[5:0];
  _RAND_39 = {1{`RANDOM}};
  replStateReg_38 = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
  replStateReg_39 = _RAND_40[5:0];
  _RAND_41 = {1{`RANDOM}};
  replStateReg_40 = _RAND_41[5:0];
  _RAND_42 = {1{`RANDOM}};
  replStateReg_41 = _RAND_42[5:0];
  _RAND_43 = {1{`RANDOM}};
  replStateReg_42 = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  replStateReg_43 = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  replStateReg_44 = _RAND_45[5:0];
  _RAND_46 = {1{`RANDOM}};
  replStateReg_45 = _RAND_46[5:0];
  _RAND_47 = {1{`RANDOM}};
  replStateReg_46 = _RAND_47[5:0];
  _RAND_48 = {1{`RANDOM}};
  replStateReg_47 = _RAND_48[5:0];
  _RAND_49 = {1{`RANDOM}};
  replStateReg_48 = _RAND_49[5:0];
  _RAND_50 = {1{`RANDOM}};
  replStateReg_49 = _RAND_50[5:0];
  _RAND_51 = {1{`RANDOM}};
  replStateReg_50 = _RAND_51[5:0];
  _RAND_52 = {1{`RANDOM}};
  replStateReg_51 = _RAND_52[5:0];
  _RAND_53 = {1{`RANDOM}};
  replStateReg_52 = _RAND_53[5:0];
  _RAND_54 = {1{`RANDOM}};
  replStateReg_53 = _RAND_54[5:0];
  _RAND_55 = {1{`RANDOM}};
  replStateReg_54 = _RAND_55[5:0];
  _RAND_56 = {1{`RANDOM}};
  replStateReg_55 = _RAND_56[5:0];
  _RAND_57 = {1{`RANDOM}};
  replStateReg_56 = _RAND_57[5:0];
  _RAND_58 = {1{`RANDOM}};
  replStateReg_57 = _RAND_58[5:0];
  _RAND_59 = {1{`RANDOM}};
  replStateReg_58 = _RAND_59[5:0];
  _RAND_60 = {1{`RANDOM}};
  replStateReg_59 = _RAND_60[5:0];
  _RAND_61 = {1{`RANDOM}};
  replStateReg_60 = _RAND_61[5:0];
  _RAND_62 = {1{`RANDOM}};
  replStateReg_61 = _RAND_62[5:0];
  _RAND_63 = {1{`RANDOM}};
  replStateReg_62 = _RAND_63[5:0];
  _RAND_64 = {1{`RANDOM}};
  replStateReg_63 = _RAND_64[5:0];
  _RAND_65 = {1{`RANDOM}};
  wayInputCache = _RAND_65[3:0];
  _RAND_66 = {1{`RANDOM}};
  tbeFields_0 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  _T_194 = _RAND_67[5:0];
  _RAND_68 = {1{`RANDOM}};
  inputToPC_addr = _RAND_68[31:0];
  _RAND_69 = {2{`RANDOM}};
  inputToPC_data = _RAND_69[63:0];
  _RAND_70 = {1{`RANDOM}};
  _T_266 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  _T_268 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  _T_269 = _RAND_72[31:0];
  _RAND_73 = {2{`RANDOM}};
  _T_270 = _RAND_73[63:0];
  _RAND_74 = {1{`RANDOM}};
  _T_273 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  _T_281 = _RAND_75[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      instUsed <= 1'h0;
    end else begin
      instUsed <= _T_83;
    end
    if (reset) begin
      replStateReg_0 <= 6'h0;
    end else if (missLD) begin
      if (6'h0 == addrReplacer[5:0]) begin
        replStateReg_0 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_1 <= 6'h0;
    end else if (missLD) begin
      if (6'h1 == addrReplacer[5:0]) begin
        replStateReg_1 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_2 <= 6'h0;
    end else if (missLD) begin
      if (6'h2 == addrReplacer[5:0]) begin
        replStateReg_2 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_3 <= 6'h0;
    end else if (missLD) begin
      if (6'h3 == addrReplacer[5:0]) begin
        replStateReg_3 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_4 <= 6'h0;
    end else if (missLD) begin
      if (6'h4 == addrReplacer[5:0]) begin
        replStateReg_4 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_5 <= 6'h0;
    end else if (missLD) begin
      if (6'h5 == addrReplacer[5:0]) begin
        replStateReg_5 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_6 <= 6'h0;
    end else if (missLD) begin
      if (6'h6 == addrReplacer[5:0]) begin
        replStateReg_6 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_7 <= 6'h0;
    end else if (missLD) begin
      if (6'h7 == addrReplacer[5:0]) begin
        replStateReg_7 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_8 <= 6'h0;
    end else if (missLD) begin
      if (6'h8 == addrReplacer[5:0]) begin
        replStateReg_8 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_9 <= 6'h0;
    end else if (missLD) begin
      if (6'h9 == addrReplacer[5:0]) begin
        replStateReg_9 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_10 <= 6'h0;
    end else if (missLD) begin
      if (6'ha == addrReplacer[5:0]) begin
        replStateReg_10 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_11 <= 6'h0;
    end else if (missLD) begin
      if (6'hb == addrReplacer[5:0]) begin
        replStateReg_11 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_12 <= 6'h0;
    end else if (missLD) begin
      if (6'hc == addrReplacer[5:0]) begin
        replStateReg_12 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_13 <= 6'h0;
    end else if (missLD) begin
      if (6'hd == addrReplacer[5:0]) begin
        replStateReg_13 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_14 <= 6'h0;
    end else if (missLD) begin
      if (6'he == addrReplacer[5:0]) begin
        replStateReg_14 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_15 <= 6'h0;
    end else if (missLD) begin
      if (6'hf == addrReplacer[5:0]) begin
        replStateReg_15 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_16 <= 6'h0;
    end else if (missLD) begin
      if (6'h10 == addrReplacer[5:0]) begin
        replStateReg_16 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_17 <= 6'h0;
    end else if (missLD) begin
      if (6'h11 == addrReplacer[5:0]) begin
        replStateReg_17 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_18 <= 6'h0;
    end else if (missLD) begin
      if (6'h12 == addrReplacer[5:0]) begin
        replStateReg_18 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_19 <= 6'h0;
    end else if (missLD) begin
      if (6'h13 == addrReplacer[5:0]) begin
        replStateReg_19 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_20 <= 6'h0;
    end else if (missLD) begin
      if (6'h14 == addrReplacer[5:0]) begin
        replStateReg_20 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_21 <= 6'h0;
    end else if (missLD) begin
      if (6'h15 == addrReplacer[5:0]) begin
        replStateReg_21 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_22 <= 6'h0;
    end else if (missLD) begin
      if (6'h16 == addrReplacer[5:0]) begin
        replStateReg_22 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_23 <= 6'h0;
    end else if (missLD) begin
      if (6'h17 == addrReplacer[5:0]) begin
        replStateReg_23 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_24 <= 6'h0;
    end else if (missLD) begin
      if (6'h18 == addrReplacer[5:0]) begin
        replStateReg_24 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_25 <= 6'h0;
    end else if (missLD) begin
      if (6'h19 == addrReplacer[5:0]) begin
        replStateReg_25 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_26 <= 6'h0;
    end else if (missLD) begin
      if (6'h1a == addrReplacer[5:0]) begin
        replStateReg_26 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_27 <= 6'h0;
    end else if (missLD) begin
      if (6'h1b == addrReplacer[5:0]) begin
        replStateReg_27 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_28 <= 6'h0;
    end else if (missLD) begin
      if (6'h1c == addrReplacer[5:0]) begin
        replStateReg_28 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_29 <= 6'h0;
    end else if (missLD) begin
      if (6'h1d == addrReplacer[5:0]) begin
        replStateReg_29 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_30 <= 6'h0;
    end else if (missLD) begin
      if (6'h1e == addrReplacer[5:0]) begin
        replStateReg_30 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_31 <= 6'h0;
    end else if (missLD) begin
      if (6'h1f == addrReplacer[5:0]) begin
        replStateReg_31 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_32 <= 6'h0;
    end else if (missLD) begin
      if (6'h20 == addrReplacer[5:0]) begin
        replStateReg_32 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_33 <= 6'h0;
    end else if (missLD) begin
      if (6'h21 == addrReplacer[5:0]) begin
        replStateReg_33 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_34 <= 6'h0;
    end else if (missLD) begin
      if (6'h22 == addrReplacer[5:0]) begin
        replStateReg_34 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_35 <= 6'h0;
    end else if (missLD) begin
      if (6'h23 == addrReplacer[5:0]) begin
        replStateReg_35 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_36 <= 6'h0;
    end else if (missLD) begin
      if (6'h24 == addrReplacer[5:0]) begin
        replStateReg_36 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_37 <= 6'h0;
    end else if (missLD) begin
      if (6'h25 == addrReplacer[5:0]) begin
        replStateReg_37 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_38 <= 6'h0;
    end else if (missLD) begin
      if (6'h26 == addrReplacer[5:0]) begin
        replStateReg_38 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_39 <= 6'h0;
    end else if (missLD) begin
      if (6'h27 == addrReplacer[5:0]) begin
        replStateReg_39 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_40 <= 6'h0;
    end else if (missLD) begin
      if (6'h28 == addrReplacer[5:0]) begin
        replStateReg_40 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_41 <= 6'h0;
    end else if (missLD) begin
      if (6'h29 == addrReplacer[5:0]) begin
        replStateReg_41 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_42 <= 6'h0;
    end else if (missLD) begin
      if (6'h2a == addrReplacer[5:0]) begin
        replStateReg_42 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_43 <= 6'h0;
    end else if (missLD) begin
      if (6'h2b == addrReplacer[5:0]) begin
        replStateReg_43 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_44 <= 6'h0;
    end else if (missLD) begin
      if (6'h2c == addrReplacer[5:0]) begin
        replStateReg_44 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_45 <= 6'h0;
    end else if (missLD) begin
      if (6'h2d == addrReplacer[5:0]) begin
        replStateReg_45 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_46 <= 6'h0;
    end else if (missLD) begin
      if (6'h2e == addrReplacer[5:0]) begin
        replStateReg_46 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_47 <= 6'h0;
    end else if (missLD) begin
      if (6'h2f == addrReplacer[5:0]) begin
        replStateReg_47 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_48 <= 6'h0;
    end else if (missLD) begin
      if (6'h30 == addrReplacer[5:0]) begin
        replStateReg_48 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_49 <= 6'h0;
    end else if (missLD) begin
      if (6'h31 == addrReplacer[5:0]) begin
        replStateReg_49 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_50 <= 6'h0;
    end else if (missLD) begin
      if (6'h32 == addrReplacer[5:0]) begin
        replStateReg_50 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_51 <= 6'h0;
    end else if (missLD) begin
      if (6'h33 == addrReplacer[5:0]) begin
        replStateReg_51 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_52 <= 6'h0;
    end else if (missLD) begin
      if (6'h34 == addrReplacer[5:0]) begin
        replStateReg_52 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_53 <= 6'h0;
    end else if (missLD) begin
      if (6'h35 == addrReplacer[5:0]) begin
        replStateReg_53 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_54 <= 6'h0;
    end else if (missLD) begin
      if (6'h36 == addrReplacer[5:0]) begin
        replStateReg_54 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_55 <= 6'h0;
    end else if (missLD) begin
      if (6'h37 == addrReplacer[5:0]) begin
        replStateReg_55 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_56 <= 6'h0;
    end else if (missLD) begin
      if (6'h38 == addrReplacer[5:0]) begin
        replStateReg_56 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_57 <= 6'h0;
    end else if (missLD) begin
      if (6'h39 == addrReplacer[5:0]) begin
        replStateReg_57 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_58 <= 6'h0;
    end else if (missLD) begin
      if (6'h3a == addrReplacer[5:0]) begin
        replStateReg_58 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_59 <= 6'h0;
    end else if (missLD) begin
      if (6'h3b == addrReplacer[5:0]) begin
        replStateReg_59 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_60 <= 6'h0;
    end else if (missLD) begin
      if (6'h3c == addrReplacer[5:0]) begin
        replStateReg_60 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_61 <= 6'h0;
    end else if (missLD) begin
      if (6'h3d == addrReplacer[5:0]) begin
        replStateReg_61 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_62 <= 6'h0;
    end else if (missLD) begin
      if (6'h3e == addrReplacer[5:0]) begin
        replStateReg_62 <= _T_186;
      end
    end
    if (reset) begin
      replStateReg_63 <= 6'h0;
    end else if (missLD) begin
      if (6'h3f == addrReplacer[5:0]) begin
        replStateReg_63 <= _T_186;
      end
    end
    if (reset) begin
      wayInputCache <= 4'h4;
    end else if (getState) begin
      if (_T_187) begin
        wayInputCache <= {{1'd0}, probeWay_io_deq_bits};
      end else begin
        wayInputCache <= tbeWay;
      end
    end
    if (reset) begin
      tbeFields_0 <= 32'h0;
    end else if (getState) begin
      tbeFields_0 <= input__io_deq_bits_tbeOut_fields_0;
    end
    if (reset) begin
      _T_194 <= 6'h4;
    end else if (getState) begin
      _T_194 <= replacerWayWire;
    end
    if (reset) begin
      inputToPC_addr <= 32'h0;
    end else if (getState) begin
      inputToPC_addr <= input__io_deq_bits_inst_addr;
    end
    if (reset) begin
      inputToPC_data <= 64'h0;
    end else if (getState) begin
      inputToPC_data <= input__io_deq_bits_inst_data;
    end
    _T_266 <= cache_io_bipassLD_in_bits_addr;
    _T_268 <= inputArbiter_io_chosen;
    _T_269 <= inputArbiter_io_out_bits_addr;
    _T_270 <= inputArbiter_io_out_bits_data;
    _T_273 <= inputArbiter_io_chosen;
    _T_281 <= tbe_io_isFull;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_267 & _T_272) begin
          $fwrite(32'h80000002,"Cache: %d req from %d Addr: %d Data: %d\n",1'h0,_T_268,_T_269,_T_270); // @[programmableCache.scala 531:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_390 & _T_272) begin
          $fwrite(32'h80000002,"Cache: %d ",1'h0); // @[programmableCache.scala 533:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_392 & _T_272) begin
          $fwrite(32'h80000002," Load hit for addr %d\n",input__io_deq_bits_inst_addr); // @[programmableCache.scala 535:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_396 & _T_272) begin
          $fwrite(32'h80000002,"addr %d is locked\n",input__io_deq_bits_inst_addr); // @[programmableCache.scala 537:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_402 & _T_272) begin
          $fwrite(32'h80000002,"TBE is full addr %d\n",input__io_deq_bits_inst_addr); // @[programmableCache.scala 539:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_410 & _T_272) begin
          $fwrite(32'h80000002,"Hit (store probably) for addr %d\n",input__io_deq_bits_inst_addr); // @[programmableCache.scala 541:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_419 & _T_272) begin
          $fwrite(32'h80000002,"miss for addr %d\n",input__io_deq_bits_inst_addr); // @[programmableCache.scala 543:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (getState & _T_272) begin
          $fwrite(32'h80000002,"Event %d Addr: %d Data: %d\n",input__io_deq_bits_inst_event,input__io_deq_bits_inst_addr,input__io_deq_bits_inst_data); // @[programmableCache.scala 549:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_16(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_inst,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_inst,
  output [63:0] io_deq_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:0]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_7_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [7:0] ram_inst [0:0]; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_7_addr; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:0]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_7_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_7_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram_addr__T_7_addr = 1'h0;
  assign ram_addr__T_7_data = ram_addr[ram_addr__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_3_data = io_enq_bits_addr;
  assign ram_addr__T_3_addr = 1'h0;
  assign ram_addr__T_3_mask = 1'h1;
  assign ram_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst__T_7_addr = 1'h0;
  assign ram_inst__T_7_data = ram_inst[ram_inst__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst__T_3_data = io_enq_bits_inst;
  assign ram_inst__T_3_addr = 1'h0;
  assign ram_inst__T_3_mask = 1'h1;
  assign ram_inst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_7_addr = 1'h0;
  assign ram_data__T_7_data = ram_data[ram_data__T_7_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = 1'h0;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst = ram_inst__T_7_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_7_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_inst[initvar] = _RAND_1[7:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_3_en & ram_addr__T_3_mask) begin
      ram_addr[ram_addr__T_3_addr] <= ram_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst__T_3_en & ram_inst__T_3_mask) begin
      ram_inst[ram_inst__T_3_addr] <= ram_inst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_4) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Queue_17(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_inst,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_inst,
  output [63:0] io_deq_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:127]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_11_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_addr__T_11_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_addr__T_3_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_addr__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_addr__T_3_en; // @[Decoupled.scala 209:16]
  reg [7:0] ram_inst [0:127]; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_11_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_inst__T_11_addr; // @[Decoupled.scala 209:16]
  wire [7:0] ram_inst__T_3_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_inst__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_inst__T_3_en; // @[Decoupled.scala 209:16]
  reg [63:0] ram_data [0:127]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_11_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_data__T_11_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire [6:0] ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [6:0] enq_ptr_value; // @[Counter.scala 29:33]
  reg [6:0] deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [6:0] _T_5 = enq_ptr_value + 7'h1; // @[Counter.scala 39:22]
  wire [6:0] _T_7 = deq_ptr_value + 7'h1; // @[Counter.scala 39:22]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  wire  _T_10 = ~full; // @[Decoupled.scala 232:19]
  assign ram_addr__T_11_addr = deq_ptr_value;
  assign ram_addr__T_11_data = ram_addr[ram_addr__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_addr__T_3_data = io_enq_bits_addr;
  assign ram_addr__T_3_addr = enq_ptr_value;
  assign ram_addr__T_3_mask = 1'h1;
  assign ram_addr__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_inst__T_11_addr = deq_ptr_value;
  assign ram_inst__T_11_data = ram_inst[ram_inst__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_inst__T_3_data = io_enq_bits_inst;
  assign ram_inst__T_3_addr = enq_ptr_value;
  assign ram_inst__T_3_mask = 1'h1;
  assign ram_inst__T_3_en = io_enq_ready & io_enq_valid;
  assign ram_data__T_11_addr = deq_ptr_value;
  assign ram_data__T_11_data = ram_data[ram_data__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = enq_ptr_value;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | _T_10; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_addr = ram_addr__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_inst = ram_inst__T_11_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = ram_data__T_11_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_inst[initvar] = _RAND_1[7:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_addr__T_3_en & ram_addr__T_3_mask) begin
      ram_addr[ram_addr__T_3_addr] <= ram_addr__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_inst__T_3_en & ram_inst__T_3_mask) begin
      ram_inst[ram_inst__T_3_addr] <= ram_inst__T_3_data; // @[Decoupled.scala 209:16]
    end
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 7'h0;
    end else if (do_enq) begin
      enq_ptr_value <= _T_5;
    end
    if (reset) begin
      deq_ptr_value <= 7'h0;
    end else if (do_deq) begin
      deq_ptr_value <= _T_7;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module CacheNode(
  input         clock,
  input         reset,
  output        io_in_cpu_ready,
  input         io_in_cpu_valid,
  input  [31:0] io_in_cpu_bits_addr,
  input  [7:0]  io_in_cpu_bits_inst,
  input  [63:0] io_in_cpu_bits_data,
  output        io_in_network_ready,
  input         io_in_network_valid,
  input  [31:0] io_in_network_bits_addr,
  input  [7:0]  io_in_network_bits_inst,
  input  [63:0] io_in_network_bits_data,
  input  [1:0]  io_in_network_bits_msgType,
  output        io_out_network_valid,
  output [31:0] io_out_network_bits_addr,
  output [7:0]  io_out_network_bits_inst,
  output [63:0] io_out_network_bits_data,
  output        io_out_cpu_valid,
  output [31:0] io_out_cpu_bits_addr,
  output        _T_297,
  output        _T_291,
  output        _T_304,
  output        hitLD,
  output        missLD,
  output        _T_294
);
  wire  cache_clock; // @[cacheNode.scala 33:21]
  wire  cache_reset; // @[cacheNode.scala 33:21]
  wire  cache_io_in_cpu_ready; // @[cacheNode.scala 33:21]
  wire  cache_io_in_cpu_valid; // @[cacheNode.scala 33:21]
  wire [1:0] cache_io_in_cpu_bits_event; // @[cacheNode.scala 33:21]
  wire [31:0] cache_io_in_cpu_bits_addr; // @[cacheNode.scala 33:21]
  wire [63:0] cache_io_in_cpu_bits_data; // @[cacheNode.scala 33:21]
  wire  cache_io_in_memCtrl_ready; // @[cacheNode.scala 33:21]
  wire  cache_io_in_memCtrl_valid; // @[cacheNode.scala 33:21]
  wire [1:0] cache_io_in_memCtrl_bits_event; // @[cacheNode.scala 33:21]
  wire [31:0] cache_io_in_memCtrl_bits_addr; // @[cacheNode.scala 33:21]
  wire [63:0] cache_io_in_memCtrl_bits_data; // @[cacheNode.scala 33:21]
  wire  cache_io_in_otherNodes_ready; // @[cacheNode.scala 33:21]
  wire  cache_io_in_otherNodes_valid; // @[cacheNode.scala 33:21]
  wire [1:0] cache_io_in_otherNodes_bits_event; // @[cacheNode.scala 33:21]
  wire [31:0] cache_io_in_otherNodes_bits_addr; // @[cacheNode.scala 33:21]
  wire [63:0] cache_io_in_otherNodes_bits_data; // @[cacheNode.scala 33:21]
  wire  cache_io_out_req_valid; // @[cacheNode.scala 33:21]
  wire [31:0] cache_io_out_req_bits_req_addr; // @[cacheNode.scala 33:21]
  wire [7:0] cache_io_out_req_bits_req_inst; // @[cacheNode.scala 33:21]
  wire [63:0] cache_io_out_req_bits_req_data; // @[cacheNode.scala 33:21]
  wire  cache_io_out_resp_valid; // @[cacheNode.scala 33:21]
  wire [31:0] cache_io_out_resp_bits_addr; // @[cacheNode.scala 33:21]
  wire  cache__T_297_0; // @[cacheNode.scala 33:21]
  wire  cache__T_291_0; // @[cacheNode.scala 33:21]
  wire  cache__T_304_0; // @[cacheNode.scala 33:21]
  wire  cache_hitLD_0; // @[cacheNode.scala 33:21]
  wire  cache_missLD_0; // @[cacheNode.scala 33:21]
  wire  cache__T_294_0; // @[cacheNode.scala 33:21]
  wire  cpuQueue_clock; // @[cacheNode.scala 34:24]
  wire  cpuQueue_reset; // @[cacheNode.scala 34:24]
  wire  cpuQueue_io_enq_ready; // @[cacheNode.scala 34:24]
  wire  cpuQueue_io_enq_valid; // @[cacheNode.scala 34:24]
  wire [31:0] cpuQueue_io_enq_bits_addr; // @[cacheNode.scala 34:24]
  wire [7:0] cpuQueue_io_enq_bits_inst; // @[cacheNode.scala 34:24]
  wire [63:0] cpuQueue_io_enq_bits_data; // @[cacheNode.scala 34:24]
  wire  cpuQueue_io_deq_ready; // @[cacheNode.scala 34:24]
  wire  cpuQueue_io_deq_valid; // @[cacheNode.scala 34:24]
  wire [31:0] cpuQueue_io_deq_bits_addr; // @[cacheNode.scala 34:24]
  wire [7:0] cpuQueue_io_deq_bits_inst; // @[cacheNode.scala 34:24]
  wire [63:0] cpuQueue_io_deq_bits_data; // @[cacheNode.scala 34:24]
  wire  memCtrlQueue_clock; // @[cacheNode.scala 35:28]
  wire  memCtrlQueue_reset; // @[cacheNode.scala 35:28]
  wire  memCtrlQueue_io_enq_ready; // @[cacheNode.scala 35:28]
  wire  memCtrlQueue_io_enq_valid; // @[cacheNode.scala 35:28]
  wire [31:0] memCtrlQueue_io_enq_bits_addr; // @[cacheNode.scala 35:28]
  wire [7:0] memCtrlQueue_io_enq_bits_inst; // @[cacheNode.scala 35:28]
  wire [63:0] memCtrlQueue_io_enq_bits_data; // @[cacheNode.scala 35:28]
  wire  memCtrlQueue_io_deq_ready; // @[cacheNode.scala 35:28]
  wire  memCtrlQueue_io_deq_valid; // @[cacheNode.scala 35:28]
  wire [31:0] memCtrlQueue_io_deq_bits_addr; // @[cacheNode.scala 35:28]
  wire [7:0] memCtrlQueue_io_deq_bits_inst; // @[cacheNode.scala 35:28]
  wire [63:0] memCtrlQueue_io_deq_bits_data; // @[cacheNode.scala 35:28]
  wire  otherNodesQueue_clock; // @[cacheNode.scala 36:31]
  wire  otherNodesQueue_reset; // @[cacheNode.scala 36:31]
  wire  otherNodesQueue_io_enq_ready; // @[cacheNode.scala 36:31]
  wire  otherNodesQueue_io_enq_valid; // @[cacheNode.scala 36:31]
  wire [31:0] otherNodesQueue_io_enq_bits_addr; // @[cacheNode.scala 36:31]
  wire [7:0] otherNodesQueue_io_enq_bits_inst; // @[cacheNode.scala 36:31]
  wire [63:0] otherNodesQueue_io_enq_bits_data; // @[cacheNode.scala 36:31]
  wire  otherNodesQueue_io_deq_ready; // @[cacheNode.scala 36:31]
  wire  otherNodesQueue_io_deq_valid; // @[cacheNode.scala 36:31]
  wire [31:0] otherNodesQueue_io_deq_bits_addr; // @[cacheNode.scala 36:31]
  wire [7:0] otherNodesQueue_io_deq_bits_inst; // @[cacheNode.scala 36:31]
  wire [63:0] otherNodesQueue_io_deq_bits_data; // @[cacheNode.scala 36:31]
  wire  _T_1 = io_in_network_ready & io_in_network_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_in_network_bits_msgType == 2'h0; // @[cacheNode.scala 54:37]
  wire  _T_3 = io_in_network_bits_msgType == 2'h1; // @[cacheNode.scala 56:43]
  wire  _GEN_2 = _T_2 ? 1'h0 : _T_3; // @[cacheNode.scala 54:45]
  programmableCache cache ( // @[cacheNode.scala 33:21]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_in_cpu_ready(cache_io_in_cpu_ready),
    .io_in_cpu_valid(cache_io_in_cpu_valid),
    .io_in_cpu_bits_event(cache_io_in_cpu_bits_event),
    .io_in_cpu_bits_addr(cache_io_in_cpu_bits_addr),
    .io_in_cpu_bits_data(cache_io_in_cpu_bits_data),
    .io_in_memCtrl_ready(cache_io_in_memCtrl_ready),
    .io_in_memCtrl_valid(cache_io_in_memCtrl_valid),
    .io_in_memCtrl_bits_event(cache_io_in_memCtrl_bits_event),
    .io_in_memCtrl_bits_addr(cache_io_in_memCtrl_bits_addr),
    .io_in_memCtrl_bits_data(cache_io_in_memCtrl_bits_data),
    .io_in_otherNodes_ready(cache_io_in_otherNodes_ready),
    .io_in_otherNodes_valid(cache_io_in_otherNodes_valid),
    .io_in_otherNodes_bits_event(cache_io_in_otherNodes_bits_event),
    .io_in_otherNodes_bits_addr(cache_io_in_otherNodes_bits_addr),
    .io_in_otherNodes_bits_data(cache_io_in_otherNodes_bits_data),
    .io_out_req_valid(cache_io_out_req_valid),
    .io_out_req_bits_req_addr(cache_io_out_req_bits_req_addr),
    .io_out_req_bits_req_inst(cache_io_out_req_bits_req_inst),
    .io_out_req_bits_req_data(cache_io_out_req_bits_req_data),
    .io_out_resp_valid(cache_io_out_resp_valid),
    .io_out_resp_bits_addr(cache_io_out_resp_bits_addr),
    ._T_297_0(cache__T_297_0),
    ._T_291_0(cache__T_291_0),
    ._T_304_0(cache__T_304_0),
    .hitLD_0(cache_hitLD_0),
    .missLD_0(cache_missLD_0),
    ._T_294_0(cache__T_294_0)
  );
  Queue_16 cpuQueue ( // @[cacheNode.scala 34:24]
    .clock(cpuQueue_clock),
    .reset(cpuQueue_reset),
    .io_enq_ready(cpuQueue_io_enq_ready),
    .io_enq_valid(cpuQueue_io_enq_valid),
    .io_enq_bits_addr(cpuQueue_io_enq_bits_addr),
    .io_enq_bits_inst(cpuQueue_io_enq_bits_inst),
    .io_enq_bits_data(cpuQueue_io_enq_bits_data),
    .io_deq_ready(cpuQueue_io_deq_ready),
    .io_deq_valid(cpuQueue_io_deq_valid),
    .io_deq_bits_addr(cpuQueue_io_deq_bits_addr),
    .io_deq_bits_inst(cpuQueue_io_deq_bits_inst),
    .io_deq_bits_data(cpuQueue_io_deq_bits_data)
  );
  Queue_17 memCtrlQueue ( // @[cacheNode.scala 35:28]
    .clock(memCtrlQueue_clock),
    .reset(memCtrlQueue_reset),
    .io_enq_ready(memCtrlQueue_io_enq_ready),
    .io_enq_valid(memCtrlQueue_io_enq_valid),
    .io_enq_bits_addr(memCtrlQueue_io_enq_bits_addr),
    .io_enq_bits_inst(memCtrlQueue_io_enq_bits_inst),
    .io_enq_bits_data(memCtrlQueue_io_enq_bits_data),
    .io_deq_ready(memCtrlQueue_io_deq_ready),
    .io_deq_valid(memCtrlQueue_io_deq_valid),
    .io_deq_bits_addr(memCtrlQueue_io_deq_bits_addr),
    .io_deq_bits_inst(memCtrlQueue_io_deq_bits_inst),
    .io_deq_bits_data(memCtrlQueue_io_deq_bits_data)
  );
  Queue_16 otherNodesQueue ( // @[cacheNode.scala 36:31]
    .clock(otherNodesQueue_clock),
    .reset(otherNodesQueue_reset),
    .io_enq_ready(otherNodesQueue_io_enq_ready),
    .io_enq_valid(otherNodesQueue_io_enq_valid),
    .io_enq_bits_addr(otherNodesQueue_io_enq_bits_addr),
    .io_enq_bits_inst(otherNodesQueue_io_enq_bits_inst),
    .io_enq_bits_data(otherNodesQueue_io_enq_bits_data),
    .io_deq_ready(otherNodesQueue_io_deq_ready),
    .io_deq_valid(otherNodesQueue_io_deq_valid),
    .io_deq_bits_addr(otherNodesQueue_io_deq_bits_addr),
    .io_deq_bits_inst(otherNodesQueue_io_deq_bits_inst),
    .io_deq_bits_data(otherNodesQueue_io_deq_bits_data)
  );
  assign io_in_cpu_ready = cpuQueue_io_enq_ready; // @[cacheNode.scala 38:19]
  assign io_in_network_ready = memCtrlQueue_io_enq_ready & otherNodesQueue_io_enq_ready; // @[cacheNode.scala 47:23]
  assign io_out_network_valid = cache_io_out_req_valid; // @[cacheNode.scala 81:24]
  assign io_out_network_bits_addr = cache_io_out_req_bits_req_addr; // @[cacheNode.scala 86:28]
  assign io_out_network_bits_inst = cache_io_out_req_bits_req_inst; // @[cacheNode.scala 84:27]
  assign io_out_network_bits_data = cache_io_out_req_bits_req_data; // @[cacheNode.scala 85:28]
  assign io_out_cpu_valid = cache_io_out_resp_valid; // @[cacheNode.scala 92:20]
  assign io_out_cpu_bits_addr = cache_io_out_resp_bits_addr; // @[cacheNode.scala 90:24]
  assign _T_297 = cache__T_297_0;
  assign _T_291 = cache__T_291_0;
  assign _T_304 = cache__T_304_0;
  assign hitLD = cache_hitLD_0;
  assign missLD = cache_missLD_0;
  assign _T_294 = cache__T_294_0;
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_in_cpu_valid = cpuQueue_io_deq_valid; // @[cacheNode.scala 64:30]
  assign cache_io_in_cpu_bits_event = cpuQueue_io_deq_bits_inst[1:0]; // @[cacheNode.scala 61:30]
  assign cache_io_in_cpu_bits_addr = cpuQueue_io_deq_bits_addr; // @[cacheNode.scala 62:30]
  assign cache_io_in_cpu_bits_data = cpuQueue_io_deq_bits_data; // @[cacheNode.scala 63:30]
  assign cache_io_in_memCtrl_valid = memCtrlQueue_io_deq_valid; // @[cacheNode.scala 70:34]
  assign cache_io_in_memCtrl_bits_event = memCtrlQueue_io_deq_bits_inst[1:0]; // @[cacheNode.scala 67:34]
  assign cache_io_in_memCtrl_bits_addr = memCtrlQueue_io_deq_bits_addr; // @[cacheNode.scala 68:34]
  assign cache_io_in_memCtrl_bits_data = memCtrlQueue_io_deq_bits_data; // @[cacheNode.scala 69:34]
  assign cache_io_in_otherNodes_valid = otherNodesQueue_io_deq_valid; // @[cacheNode.scala 76:37]
  assign cache_io_in_otherNodes_bits_event = otherNodesQueue_io_deq_bits_inst[1:0]; // @[cacheNode.scala 73:37]
  assign cache_io_in_otherNodes_bits_addr = otherNodesQueue_io_deq_bits_addr; // @[cacheNode.scala 74:37]
  assign cache_io_in_otherNodes_bits_data = otherNodesQueue_io_deq_bits_data; // @[cacheNode.scala 75:37]
  assign cpuQueue_clock = clock;
  assign cpuQueue_reset = reset;
  assign cpuQueue_io_enq_valid = io_in_cpu_valid; // @[cacheNode.scala 38:19]
  assign cpuQueue_io_enq_bits_addr = io_in_cpu_bits_addr; // @[cacheNode.scala 38:19]
  assign cpuQueue_io_enq_bits_inst = io_in_cpu_bits_inst; // @[cacheNode.scala 38:19]
  assign cpuQueue_io_enq_bits_data = io_in_cpu_bits_data; // @[cacheNode.scala 38:19]
  assign cpuQueue_io_deq_ready = cache_io_in_cpu_ready; // @[cacheNode.scala 65:25]
  assign memCtrlQueue_clock = clock;
  assign memCtrlQueue_reset = reset;
  assign memCtrlQueue_io_enq_valid = _T_1 & _T_2; // @[cacheNode.scala 49:29 cacheNode.scala 55:33]
  assign memCtrlQueue_io_enq_bits_addr = io_in_network_bits_addr; // @[cacheNode.scala 39:33]
  assign memCtrlQueue_io_enq_bits_inst = io_in_network_bits_inst; // @[cacheNode.scala 41:33]
  assign memCtrlQueue_io_enq_bits_data = io_in_network_bits_data; // @[cacheNode.scala 40:33]
  assign memCtrlQueue_io_deq_ready = cache_io_in_memCtrl_ready; // @[cacheNode.scala 71:29]
  assign otherNodesQueue_clock = clock;
  assign otherNodesQueue_reset = reset;
  assign otherNodesQueue_io_enq_valid = _T_1 & _GEN_2; // @[cacheNode.scala 50:32 cacheNode.scala 57:36]
  assign otherNodesQueue_io_enq_bits_addr = io_in_network_bits_addr; // @[cacheNode.scala 43:36]
  assign otherNodesQueue_io_enq_bits_inst = io_in_network_bits_inst; // @[cacheNode.scala 45:36]
  assign otherNodesQueue_io_enq_bits_data = io_in_network_bits_data; // @[cacheNode.scala 44:36]
  assign otherNodesQueue_io_deq_ready = cache_io_in_otherNodes_ready; // @[cacheNode.scala 77:32]
endmodule
module Bore(
  input         clock,
  input         reset,
  output [31:0] io_events_0,
  output [31:0] io_events_1,
  output [31:0] io_events_2,
  output [31:0] io_events_3,
  output [31:0] io_events_4,
  output [31:0] io_events_5,
  input         memCtrlReq_0,
  input         instCount_0,
  input         ldReq_0,
  input         hitLD_0,
  input         missLD_0,
  input         cpuReq_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [23:0] _T_1; // @[Counter.scala 29:33]
  wire  _T_3 = _T_1 == 24'h98967f; // @[Counter.scala 38:24]
  wire [23:0] _T_5 = _T_1 + 24'h1; // @[Counter.scala 39:22]
  reg [23:0] _T_6; // @[Counter.scala 29:33]
  wire  _T_8 = _T_6 == 24'h98967f; // @[Counter.scala 38:24]
  wire [23:0] _T_10 = _T_6 + 24'h1; // @[Counter.scala 39:22]
  reg [23:0] _T_11; // @[Counter.scala 29:33]
  wire  _T_13 = _T_11 == 24'h98967f; // @[Counter.scala 38:24]
  wire [23:0] _T_15 = _T_11 + 24'h1; // @[Counter.scala 39:22]
  reg [23:0] _T_16; // @[Counter.scala 29:33]
  wire  _T_18 = _T_16 == 24'h98967f; // @[Counter.scala 38:24]
  wire [23:0] _T_20 = _T_16 + 24'h1; // @[Counter.scala 39:22]
  reg [23:0] _T_21; // @[Counter.scala 29:33]
  wire  _T_23 = _T_21 == 24'h98967f; // @[Counter.scala 38:24]
  wire [23:0] _T_25 = _T_21 + 24'h1; // @[Counter.scala 39:22]
  reg [23:0] _T_26; // @[Counter.scala 29:33]
  wire  _T_28 = _T_26 == 24'h98967f; // @[Counter.scala 38:24]
  wire [23:0] _T_30 = _T_26 + 24'h1; // @[Counter.scala 39:22]
  assign io_events_0 = {{8'd0}, _T_1}; // @[memGenTopLevel.scala 40:15]
  assign io_events_1 = {{8'd0}, _T_6}; // @[memGenTopLevel.scala 40:15]
  assign io_events_2 = {{8'd0}, _T_11}; // @[memGenTopLevel.scala 40:15]
  assign io_events_3 = {{8'd0}, _T_16}; // @[memGenTopLevel.scala 40:15]
  assign io_events_4 = {{8'd0}, _T_21}; // @[memGenTopLevel.scala 40:15]
  assign io_events_5 = {{8'd0}, _T_26}; // @[memGenTopLevel.scala 40:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[23:0];
  _RAND_1 = {1{`RANDOM}};
  _T_6 = _RAND_1[23:0];
  _RAND_2 = {1{`RANDOM}};
  _T_11 = _RAND_2[23:0];
  _RAND_3 = {1{`RANDOM}};
  _T_16 = _RAND_3[23:0];
  _RAND_4 = {1{`RANDOM}};
  _T_21 = _RAND_4[23:0];
  _RAND_5 = {1{`RANDOM}};
  _T_26 = _RAND_5[23:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1 <= 24'h0;
    end else if (missLD_0) begin
      if (_T_3) begin
        _T_1 <= 24'h0;
      end else begin
        _T_1 <= _T_5;
      end
    end
    if (reset) begin
      _T_6 <= 24'h0;
    end else if (hitLD_0) begin
      if (_T_8) begin
        _T_6 <= 24'h0;
      end else begin
        _T_6 <= _T_10;
      end
    end
    if (reset) begin
      _T_11 <= 24'h0;
    end else if (instCount_0) begin
      if (_T_13) begin
        _T_11 <= 24'h0;
      end else begin
        _T_11 <= _T_15;
      end
    end
    if (reset) begin
      _T_16 <= 24'h0;
    end else if (cpuReq_0) begin
      if (_T_18) begin
        _T_16 <= 24'h0;
      end else begin
        _T_16 <= _T_20;
      end
    end
    if (reset) begin
      _T_21 <= 24'h0;
    end else if (memCtrlReq_0) begin
      if (_T_23) begin
        _T_21 <= 24'h0;
      end else begin
        _T_21 <= _T_25;
      end
    end
    if (reset) begin
      _T_26 <= 24'h0;
    end else if (ldReq_0) begin
      if (_T_28) begin
        _T_26 <= 24'h0;
      end else begin
        _T_26 <= _T_30;
      end
    end
  end
endmodule
module memGenTopLevel(
  input         clock,
  input         reset,
  output        io_instruction_0_ready,
  input         io_instruction_0_valid,
  input  [31:0] io_instruction_0_bits_addr,
  input  [7:0]  io_instruction_0_bits_inst,
  input  [63:0] io_instruction_0_bits_data,
  output        io_resp_0_valid,
  output [31:0] io_resp_0_bits_addr,
  output [31:0] io_events_bits_0,
  output [31:0] io_events_bits_1,
  output [31:0] io_events_bits_2,
  output [31:0] io_events_bits_3,
  output [31:0] io_events_bits_4,
  output [31:0] io_events_bits_5,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output        io_mem_b_ready,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [15:0] io_mem_ar_bits_len,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last
);
  wire  memCtrl_clock; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_reset; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_in_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_in_valid; // @[memGenTopLevel.scala 67:25]
  wire [31:0] memCtrl_io_in_bits_addr; // @[memGenTopLevel.scala 67:25]
  wire [7:0] memCtrl_io_in_bits_inst; // @[memGenTopLevel.scala 67:25]
  wire [63:0] memCtrl_io_in_bits_data; // @[memGenTopLevel.scala 67:25]
  wire [2:0] memCtrl_io_in_bits_src; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_aw_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_aw_valid; // @[memGenTopLevel.scala 67:25]
  wire [31:0] memCtrl_io_mem_aw_bits_addr; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_w_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_w_valid; // @[memGenTopLevel.scala 67:25]
  wire [63:0] memCtrl_io_mem_w_bits_data; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_b_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_ar_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_ar_valid; // @[memGenTopLevel.scala 67:25]
  wire [31:0] memCtrl_io_mem_ar_bits_addr; // @[memGenTopLevel.scala 67:25]
  wire [15:0] memCtrl_io_mem_ar_bits_len; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_r_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_r_valid; // @[memGenTopLevel.scala 67:25]
  wire [63:0] memCtrl_io_mem_r_bits_data; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_mem_r_bits_last; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_out_ready; // @[memGenTopLevel.scala 67:25]
  wire  memCtrl_io_out_valid; // @[memGenTopLevel.scala 67:25]
  wire [31:0] memCtrl_io_out_bits_addr; // @[memGenTopLevel.scala 67:25]
  wire [63:0] memCtrl_io_out_bits_data; // @[memGenTopLevel.scala 67:25]
  wire [2:0] memCtrl_io_out_bits_dst; // @[memGenTopLevel.scala 67:25]
  wire  memCtrlInputQueue_clock; // @[memGenTopLevel.scala 68:35]
  wire  memCtrlInputQueue_reset; // @[memGenTopLevel.scala 68:35]
  wire  memCtrlInputQueue_io_enq_ready; // @[memGenTopLevel.scala 68:35]
  wire  memCtrlInputQueue_io_enq_valid; // @[memGenTopLevel.scala 68:35]
  wire [31:0] memCtrlInputQueue_io_enq_bits_addr; // @[memGenTopLevel.scala 68:35]
  wire [7:0] memCtrlInputQueue_io_enq_bits_inst; // @[memGenTopLevel.scala 68:35]
  wire [63:0] memCtrlInputQueue_io_enq_bits_data; // @[memGenTopLevel.scala 68:35]
  wire [2:0] memCtrlInputQueue_io_enq_bits_src; // @[memGenTopLevel.scala 68:35]
  wire  memCtrlInputQueue_io_deq_ready; // @[memGenTopLevel.scala 68:35]
  wire  memCtrlInputQueue_io_deq_valid; // @[memGenTopLevel.scala 68:35]
  wire [31:0] memCtrlInputQueue_io_deq_bits_addr; // @[memGenTopLevel.scala 68:35]
  wire [7:0] memCtrlInputQueue_io_deq_bits_inst; // @[memGenTopLevel.scala 68:35]
  wire [63:0] memCtrlInputQueue_io_deq_bits_data; // @[memGenTopLevel.scala 68:35]
  wire [2:0] memCtrlInputQueue_io_deq_bits_src; // @[memGenTopLevel.scala 68:35]
  wire  routerNode_0_clock; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_reset; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_cacheIn_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_0_io_cacheIn_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_0_io_cacheIn_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_0_io_cacheIn_bits_data; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_cacheOut_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_cacheOut_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_0_io_cacheOut_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_0_io_cacheOut_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_0_io_cacheOut_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [1:0] routerNode_0_io_cacheOut_bits_msgType; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_in_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_in_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_0_io_in_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_0_io_in_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_0_io_in_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_0_io_in_bits_src; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_0_io_in_bits_dst; // @[memGenTopLevel.scala 70:28]
  wire [1:0] routerNode_0_io_in_bits_msgType; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_out_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_0_io_out_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_0_io_out_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_0_io_out_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_0_io_out_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_0_io_out_bits_src; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_0_io_out_bits_dst; // @[memGenTopLevel.scala 70:28]
  wire [1:0] routerNode_0_io_out_bits_msgType; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_clock; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_reset; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_cacheIn_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_cacheIn_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_1_io_cacheIn_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_1_io_cacheIn_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_1_io_cacheIn_bits_dst; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_cacheOut_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_cacheOut_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_1_io_cacheOut_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_1_io_cacheOut_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_1_io_cacheOut_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_1_io_cacheOut_bits_src; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_in_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_in_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_1_io_in_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_1_io_in_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_1_io_in_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_1_io_in_bits_src; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_1_io_in_bits_dst; // @[memGenTopLevel.scala 70:28]
  wire [1:0] routerNode_1_io_in_bits_msgType; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_out_ready; // @[memGenTopLevel.scala 70:28]
  wire  routerNode_1_io_out_valid; // @[memGenTopLevel.scala 70:28]
  wire [31:0] routerNode_1_io_out_bits_addr; // @[memGenTopLevel.scala 70:28]
  wire [7:0] routerNode_1_io_out_bits_inst; // @[memGenTopLevel.scala 70:28]
  wire [63:0] routerNode_1_io_out_bits_data; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_1_io_out_bits_src; // @[memGenTopLevel.scala 70:28]
  wire [2:0] routerNode_1_io_out_bits_dst; // @[memGenTopLevel.scala 70:28]
  wire [1:0] routerNode_1_io_out_bits_msgType; // @[memGenTopLevel.scala 70:28]
  wire  cacheNode_0_clock; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_reset; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_io_in_cpu_ready; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_io_in_cpu_valid; // @[memGenTopLevel.scala 74:28]
  wire [31:0] cacheNode_0_io_in_cpu_bits_addr; // @[memGenTopLevel.scala 74:28]
  wire [7:0] cacheNode_0_io_in_cpu_bits_inst; // @[memGenTopLevel.scala 74:28]
  wire [63:0] cacheNode_0_io_in_cpu_bits_data; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_io_in_network_ready; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_io_in_network_valid; // @[memGenTopLevel.scala 74:28]
  wire [31:0] cacheNode_0_io_in_network_bits_addr; // @[memGenTopLevel.scala 74:28]
  wire [7:0] cacheNode_0_io_in_network_bits_inst; // @[memGenTopLevel.scala 74:28]
  wire [63:0] cacheNode_0_io_in_network_bits_data; // @[memGenTopLevel.scala 74:28]
  wire [1:0] cacheNode_0_io_in_network_bits_msgType; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_io_out_network_valid; // @[memGenTopLevel.scala 74:28]
  wire [31:0] cacheNode_0_io_out_network_bits_addr; // @[memGenTopLevel.scala 74:28]
  wire [7:0] cacheNode_0_io_out_network_bits_inst; // @[memGenTopLevel.scala 74:28]
  wire [63:0] cacheNode_0_io_out_network_bits_data; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_io_out_cpu_valid; // @[memGenTopLevel.scala 74:28]
  wire [31:0] cacheNode_0_io_out_cpu_bits_addr; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0__T_297; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0__T_291; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0__T_304; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_hitLD; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0_missLD; // @[memGenTopLevel.scala 74:28]
  wire  cacheNode_0__T_294; // @[memGenTopLevel.scala 74:28]
  wire  bore_clock; // @[memGenTopLevel.scala 78:22]
  wire  bore_reset; // @[memGenTopLevel.scala 78:22]
  wire [31:0] bore_io_events_0; // @[memGenTopLevel.scala 78:22]
  wire [31:0] bore_io_events_1; // @[memGenTopLevel.scala 78:22]
  wire [31:0] bore_io_events_2; // @[memGenTopLevel.scala 78:22]
  wire [31:0] bore_io_events_3; // @[memGenTopLevel.scala 78:22]
  wire [31:0] bore_io_events_4; // @[memGenTopLevel.scala 78:22]
  wire [31:0] bore_io_events_5; // @[memGenTopLevel.scala 78:22]
  wire  bore_memCtrlReq_0; // @[memGenTopLevel.scala 78:22]
  wire  bore_instCount_0; // @[memGenTopLevel.scala 78:22]
  wire  bore_ldReq_0; // @[memGenTopLevel.scala 78:22]
  wire  bore_hitLD_0; // @[memGenTopLevel.scala 78:22]
  wire  bore_missLD_0; // @[memGenTopLevel.scala 78:22]
  wire  bore_cpuReq_0; // @[memGenTopLevel.scala 78:22]
  memoryWrapper memCtrl ( // @[memGenTopLevel.scala 67:25]
    .clock(memCtrl_clock),
    .reset(memCtrl_reset),
    .io_in_ready(memCtrl_io_in_ready),
    .io_in_valid(memCtrl_io_in_valid),
    .io_in_bits_addr(memCtrl_io_in_bits_addr),
    .io_in_bits_inst(memCtrl_io_in_bits_inst),
    .io_in_bits_data(memCtrl_io_in_bits_data),
    .io_in_bits_src(memCtrl_io_in_bits_src),
    .io_mem_aw_ready(memCtrl_io_mem_aw_ready),
    .io_mem_aw_valid(memCtrl_io_mem_aw_valid),
    .io_mem_aw_bits_addr(memCtrl_io_mem_aw_bits_addr),
    .io_mem_w_ready(memCtrl_io_mem_w_ready),
    .io_mem_w_valid(memCtrl_io_mem_w_valid),
    .io_mem_w_bits_data(memCtrl_io_mem_w_bits_data),
    .io_mem_b_ready(memCtrl_io_mem_b_ready),
    .io_mem_ar_ready(memCtrl_io_mem_ar_ready),
    .io_mem_ar_valid(memCtrl_io_mem_ar_valid),
    .io_mem_ar_bits_addr(memCtrl_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(memCtrl_io_mem_ar_bits_len),
    .io_mem_r_ready(memCtrl_io_mem_r_ready),
    .io_mem_r_valid(memCtrl_io_mem_r_valid),
    .io_mem_r_bits_data(memCtrl_io_mem_r_bits_data),
    .io_mem_r_bits_last(memCtrl_io_mem_r_bits_last),
    .io_out_ready(memCtrl_io_out_ready),
    .io_out_valid(memCtrl_io_out_valid),
    .io_out_bits_addr(memCtrl_io_out_bits_addr),
    .io_out_bits_data(memCtrl_io_out_bits_data),
    .io_out_bits_dst(memCtrl_io_out_bits_dst)
  );
  Queue memCtrlInputQueue ( // @[memGenTopLevel.scala 68:35]
    .clock(memCtrlInputQueue_clock),
    .reset(memCtrlInputQueue_reset),
    .io_enq_ready(memCtrlInputQueue_io_enq_ready),
    .io_enq_valid(memCtrlInputQueue_io_enq_valid),
    .io_enq_bits_addr(memCtrlInputQueue_io_enq_bits_addr),
    .io_enq_bits_inst(memCtrlInputQueue_io_enq_bits_inst),
    .io_enq_bits_data(memCtrlInputQueue_io_enq_bits_data),
    .io_enq_bits_src(memCtrlInputQueue_io_enq_bits_src),
    .io_deq_ready(memCtrlInputQueue_io_deq_ready),
    .io_deq_valid(memCtrlInputQueue_io_deq_valid),
    .io_deq_bits_addr(memCtrlInputQueue_io_deq_bits_addr),
    .io_deq_bits_inst(memCtrlInputQueue_io_deq_bits_inst),
    .io_deq_bits_data(memCtrlInputQueue_io_deq_bits_data),
    .io_deq_bits_src(memCtrlInputQueue_io_deq_bits_src)
  );
  Router routerNode_0 ( // @[memGenTopLevel.scala 70:28]
    .clock(routerNode_0_clock),
    .reset(routerNode_0_reset),
    .io_cacheIn_valid(routerNode_0_io_cacheIn_valid),
    .io_cacheIn_bits_addr(routerNode_0_io_cacheIn_bits_addr),
    .io_cacheIn_bits_inst(routerNode_0_io_cacheIn_bits_inst),
    .io_cacheIn_bits_data(routerNode_0_io_cacheIn_bits_data),
    .io_cacheOut_ready(routerNode_0_io_cacheOut_ready),
    .io_cacheOut_valid(routerNode_0_io_cacheOut_valid),
    .io_cacheOut_bits_addr(routerNode_0_io_cacheOut_bits_addr),
    .io_cacheOut_bits_inst(routerNode_0_io_cacheOut_bits_inst),
    .io_cacheOut_bits_data(routerNode_0_io_cacheOut_bits_data),
    .io_cacheOut_bits_msgType(routerNode_0_io_cacheOut_bits_msgType),
    .io_in_ready(routerNode_0_io_in_ready),
    .io_in_valid(routerNode_0_io_in_valid),
    .io_in_bits_addr(routerNode_0_io_in_bits_addr),
    .io_in_bits_inst(routerNode_0_io_in_bits_inst),
    .io_in_bits_data(routerNode_0_io_in_bits_data),
    .io_in_bits_src(routerNode_0_io_in_bits_src),
    .io_in_bits_dst(routerNode_0_io_in_bits_dst),
    .io_in_bits_msgType(routerNode_0_io_in_bits_msgType),
    .io_out_ready(routerNode_0_io_out_ready),
    .io_out_valid(routerNode_0_io_out_valid),
    .io_out_bits_addr(routerNode_0_io_out_bits_addr),
    .io_out_bits_inst(routerNode_0_io_out_bits_inst),
    .io_out_bits_data(routerNode_0_io_out_bits_data),
    .io_out_bits_src(routerNode_0_io_out_bits_src),
    .io_out_bits_dst(routerNode_0_io_out_bits_dst),
    .io_out_bits_msgType(routerNode_0_io_out_bits_msgType)
  );
  Router_1 routerNode_1 ( // @[memGenTopLevel.scala 70:28]
    .clock(routerNode_1_clock),
    .reset(routerNode_1_reset),
    .io_cacheIn_ready(routerNode_1_io_cacheIn_ready),
    .io_cacheIn_valid(routerNode_1_io_cacheIn_valid),
    .io_cacheIn_bits_addr(routerNode_1_io_cacheIn_bits_addr),
    .io_cacheIn_bits_data(routerNode_1_io_cacheIn_bits_data),
    .io_cacheIn_bits_dst(routerNode_1_io_cacheIn_bits_dst),
    .io_cacheOut_ready(routerNode_1_io_cacheOut_ready),
    .io_cacheOut_valid(routerNode_1_io_cacheOut_valid),
    .io_cacheOut_bits_addr(routerNode_1_io_cacheOut_bits_addr),
    .io_cacheOut_bits_inst(routerNode_1_io_cacheOut_bits_inst),
    .io_cacheOut_bits_data(routerNode_1_io_cacheOut_bits_data),
    .io_cacheOut_bits_src(routerNode_1_io_cacheOut_bits_src),
    .io_in_ready(routerNode_1_io_in_ready),
    .io_in_valid(routerNode_1_io_in_valid),
    .io_in_bits_addr(routerNode_1_io_in_bits_addr),
    .io_in_bits_inst(routerNode_1_io_in_bits_inst),
    .io_in_bits_data(routerNode_1_io_in_bits_data),
    .io_in_bits_src(routerNode_1_io_in_bits_src),
    .io_in_bits_dst(routerNode_1_io_in_bits_dst),
    .io_in_bits_msgType(routerNode_1_io_in_bits_msgType),
    .io_out_ready(routerNode_1_io_out_ready),
    .io_out_valid(routerNode_1_io_out_valid),
    .io_out_bits_addr(routerNode_1_io_out_bits_addr),
    .io_out_bits_inst(routerNode_1_io_out_bits_inst),
    .io_out_bits_data(routerNode_1_io_out_bits_data),
    .io_out_bits_src(routerNode_1_io_out_bits_src),
    .io_out_bits_dst(routerNode_1_io_out_bits_dst),
    .io_out_bits_msgType(routerNode_1_io_out_bits_msgType)
  );
  CacheNode cacheNode_0 ( // @[memGenTopLevel.scala 74:28]
    .clock(cacheNode_0_clock),
    .reset(cacheNode_0_reset),
    .io_in_cpu_ready(cacheNode_0_io_in_cpu_ready),
    .io_in_cpu_valid(cacheNode_0_io_in_cpu_valid),
    .io_in_cpu_bits_addr(cacheNode_0_io_in_cpu_bits_addr),
    .io_in_cpu_bits_inst(cacheNode_0_io_in_cpu_bits_inst),
    .io_in_cpu_bits_data(cacheNode_0_io_in_cpu_bits_data),
    .io_in_network_ready(cacheNode_0_io_in_network_ready),
    .io_in_network_valid(cacheNode_0_io_in_network_valid),
    .io_in_network_bits_addr(cacheNode_0_io_in_network_bits_addr),
    .io_in_network_bits_inst(cacheNode_0_io_in_network_bits_inst),
    .io_in_network_bits_data(cacheNode_0_io_in_network_bits_data),
    .io_in_network_bits_msgType(cacheNode_0_io_in_network_bits_msgType),
    .io_out_network_valid(cacheNode_0_io_out_network_valid),
    .io_out_network_bits_addr(cacheNode_0_io_out_network_bits_addr),
    .io_out_network_bits_inst(cacheNode_0_io_out_network_bits_inst),
    .io_out_network_bits_data(cacheNode_0_io_out_network_bits_data),
    .io_out_cpu_valid(cacheNode_0_io_out_cpu_valid),
    .io_out_cpu_bits_addr(cacheNode_0_io_out_cpu_bits_addr),
    ._T_297(cacheNode_0__T_297),
    ._T_291(cacheNode_0__T_291),
    ._T_304(cacheNode_0__T_304),
    .hitLD(cacheNode_0_hitLD),
    .missLD(cacheNode_0_missLD),
    ._T_294(cacheNode_0__T_294)
  );
  Bore bore ( // @[memGenTopLevel.scala 78:22]
    .clock(bore_clock),
    .reset(bore_reset),
    .io_events_0(bore_io_events_0),
    .io_events_1(bore_io_events_1),
    .io_events_2(bore_io_events_2),
    .io_events_3(bore_io_events_3),
    .io_events_4(bore_io_events_4),
    .io_events_5(bore_io_events_5),
    .memCtrlReq_0(bore_memCtrlReq_0),
    .instCount_0(bore_instCount_0),
    .ldReq_0(bore_ldReq_0),
    .hitLD_0(bore_hitLD_0),
    .missLD_0(bore_missLD_0),
    .cpuReq_0(bore_cpuReq_0)
  );
  assign io_instruction_0_ready = cacheNode_0_io_in_cpu_ready; // @[memGenTopLevel.scala 88:33]
  assign io_resp_0_valid = cacheNode_0_io_out_cpu_valid; // @[memGenTopLevel.scala 89:20]
  assign io_resp_0_bits_addr = cacheNode_0_io_out_cpu_bits_addr; // @[memGenTopLevel.scala 89:20]
  assign io_events_bits_0 = bore_io_events_0; // @[memGenTopLevel.scala 82:20]
  assign io_events_bits_1 = bore_io_events_1; // @[memGenTopLevel.scala 82:20]
  assign io_events_bits_2 = bore_io_events_2; // @[memGenTopLevel.scala 82:20]
  assign io_events_bits_3 = bore_io_events_3; // @[memGenTopLevel.scala 82:20]
  assign io_events_bits_4 = bore_io_events_4; // @[memGenTopLevel.scala 82:20]
  assign io_events_bits_5 = bore_io_events_5; // @[memGenTopLevel.scala 82:20]
  assign io_mem_aw_valid = memCtrl_io_mem_aw_valid; // @[memGenTopLevel.scala 100:12]
  assign io_mem_aw_bits_addr = memCtrl_io_mem_aw_bits_addr; // @[memGenTopLevel.scala 100:12]
  assign io_mem_w_valid = memCtrl_io_mem_w_valid; // @[memGenTopLevel.scala 100:12]
  assign io_mem_w_bits_data = memCtrl_io_mem_w_bits_data; // @[memGenTopLevel.scala 100:12]
  assign io_mem_b_ready = memCtrl_io_mem_b_ready; // @[memGenTopLevel.scala 100:12]
  assign io_mem_ar_valid = memCtrl_io_mem_ar_valid; // @[memGenTopLevel.scala 100:12]
  assign io_mem_ar_bits_addr = memCtrl_io_mem_ar_bits_addr; // @[memGenTopLevel.scala 100:12]
  assign io_mem_ar_bits_len = memCtrl_io_mem_ar_bits_len; // @[memGenTopLevel.scala 100:12]
  assign io_mem_r_ready = memCtrl_io_mem_r_ready; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_clock = clock;
  assign memCtrl_reset = reset;
  assign memCtrl_io_in_valid = memCtrlInputQueue_io_deq_valid; // @[memGenTopLevel.scala 98:19]
  assign memCtrl_io_in_bits_addr = memCtrlInputQueue_io_deq_bits_addr; // @[memGenTopLevel.scala 98:19]
  assign memCtrl_io_in_bits_inst = memCtrlInputQueue_io_deq_bits_inst; // @[memGenTopLevel.scala 98:19]
  assign memCtrl_io_in_bits_data = memCtrlInputQueue_io_deq_bits_data; // @[memGenTopLevel.scala 98:19]
  assign memCtrl_io_in_bits_src = memCtrlInputQueue_io_deq_bits_src; // @[memGenTopLevel.scala 98:19]
  assign memCtrl_io_mem_aw_ready = io_mem_aw_ready; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_io_mem_w_ready = io_mem_w_ready; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_io_mem_ar_ready = io_mem_ar_ready; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_io_mem_r_valid = io_mem_r_valid; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_io_mem_r_bits_data = io_mem_r_bits_data; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_io_mem_r_bits_last = io_mem_r_bits_last; // @[memGenTopLevel.scala 100:12]
  assign memCtrl_io_out_ready = routerNode_1_io_cacheIn_ready; // @[memGenTopLevel.scala 99:52]
  assign memCtrlInputQueue_clock = clock;
  assign memCtrlInputQueue_reset = reset;
  assign memCtrlInputQueue_io_enq_valid = routerNode_1_io_cacheOut_valid; // @[memGenTopLevel.scala 97:30]
  assign memCtrlInputQueue_io_enq_bits_addr = routerNode_1_io_cacheOut_bits_addr; // @[memGenTopLevel.scala 97:30]
  assign memCtrlInputQueue_io_enq_bits_inst = routerNode_1_io_cacheOut_bits_inst; // @[memGenTopLevel.scala 97:30]
  assign memCtrlInputQueue_io_enq_bits_data = routerNode_1_io_cacheOut_bits_data; // @[memGenTopLevel.scala 97:30]
  assign memCtrlInputQueue_io_enq_bits_src = routerNode_1_io_cacheOut_bits_src; // @[memGenTopLevel.scala 97:30]
  assign memCtrlInputQueue_io_deq_ready = memCtrl_io_in_ready; // @[memGenTopLevel.scala 98:19]
  assign routerNode_0_clock = clock;
  assign routerNode_0_reset = reset;
  assign routerNode_0_io_cacheIn_valid = cacheNode_0_io_out_network_valid; // @[memGenTopLevel.scala 93:34]
  assign routerNode_0_io_cacheIn_bits_addr = cacheNode_0_io_out_network_bits_addr; // @[memGenTopLevel.scala 93:34]
  assign routerNode_0_io_cacheIn_bits_inst = cacheNode_0_io_out_network_bits_inst; // @[memGenTopLevel.scala 93:34]
  assign routerNode_0_io_cacheIn_bits_data = cacheNode_0_io_out_network_bits_data; // @[memGenTopLevel.scala 93:34]
  assign routerNode_0_io_cacheOut_ready = cacheNode_0_io_in_network_ready; // @[memGenTopLevel.scala 94:36]
  assign routerNode_0_io_in_valid = routerNode_1_io_out_valid; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_in_bits_addr = routerNode_1_io_out_bits_addr; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_in_bits_inst = routerNode_1_io_out_bits_inst; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_in_bits_data = routerNode_1_io_out_bits_data; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_in_bits_src = routerNode_1_io_out_bits_src; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_in_bits_dst = routerNode_1_io_out_bits_dst; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_in_bits_msgType = routerNode_1_io_out_bits_msgType; // @[memGenTopLevel.scala 105:25]
  assign routerNode_0_io_out_ready = routerNode_1_io_in_ready; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_clock = clock;
  assign routerNode_1_reset = reset;
  assign routerNode_1_io_cacheIn_valid = memCtrl_io_out_valid; // @[memGenTopLevel.scala 99:52]
  assign routerNode_1_io_cacheIn_bits_addr = memCtrl_io_out_bits_addr; // @[memGenTopLevel.scala 99:52]
  assign routerNode_1_io_cacheIn_bits_data = memCtrl_io_out_bits_data; // @[memGenTopLevel.scala 99:52]
  assign routerNode_1_io_cacheIn_bits_dst = memCtrl_io_out_bits_dst; // @[memGenTopLevel.scala 99:52]
  assign routerNode_1_io_cacheOut_ready = memCtrlInputQueue_io_enq_ready; // @[memGenTopLevel.scala 97:30]
  assign routerNode_1_io_in_valid = routerNode_0_io_out_valid; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_in_bits_addr = routerNode_0_io_out_bits_addr; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_in_bits_inst = routerNode_0_io_out_bits_inst; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_in_bits_data = routerNode_0_io_out_bits_data; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_in_bits_src = routerNode_0_io_out_bits_src; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_in_bits_dst = routerNode_0_io_out_bits_dst; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_in_bits_msgType = routerNode_0_io_out_bits_msgType; // @[memGenTopLevel.scala 103:32]
  assign routerNode_1_io_out_ready = routerNode_0_io_in_ready; // @[memGenTopLevel.scala 105:25]
  assign cacheNode_0_clock = clock;
  assign cacheNode_0_reset = reset;
  assign cacheNode_0_io_in_cpu_valid = io_instruction_0_valid; // @[memGenTopLevel.scala 87:38]
  assign cacheNode_0_io_in_cpu_bits_addr = io_instruction_0_bits_addr; // @[memGenTopLevel.scala 86:34]
  assign cacheNode_0_io_in_cpu_bits_inst = io_instruction_0_bits_inst; // @[memGenTopLevel.scala 86:34]
  assign cacheNode_0_io_in_cpu_bits_data = io_instruction_0_bits_data; // @[memGenTopLevel.scala 86:34]
  assign cacheNode_0_io_in_network_valid = routerNode_0_io_cacheOut_valid; // @[memGenTopLevel.scala 94:36]
  assign cacheNode_0_io_in_network_bits_addr = routerNode_0_io_cacheOut_bits_addr; // @[memGenTopLevel.scala 94:36]
  assign cacheNode_0_io_in_network_bits_inst = routerNode_0_io_cacheOut_bits_inst; // @[memGenTopLevel.scala 94:36]
  assign cacheNode_0_io_in_network_bits_data = routerNode_0_io_cacheOut_bits_data; // @[memGenTopLevel.scala 94:36]
  assign cacheNode_0_io_in_network_bits_msgType = routerNode_0_io_cacheOut_bits_msgType; // @[memGenTopLevel.scala 94:36]
  assign bore_clock = clock;
  assign bore_reset = reset;
  assign bore_memCtrlReq_0 = cacheNode_0__T_297;
  assign bore_instCount_0 = cacheNode_0__T_291;
  assign bore_ldReq_0 = cacheNode_0__T_304;
  assign bore_hitLD_0 = cacheNode_0_hitLD;
  assign bore_missLD_0 = cacheNode_0_missLD;
  assign bore_cpuReq_0 = cacheNode_0__T_294;
endmodule
module Arbiter_6(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits = io_in_0_bits; // @[Arbiter.scala 124:15]
endmodule
module Queue_19(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram [0:15]; // @[Decoupled.scala 209:16]
  wire [31:0] ram__T_11_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram__T_11_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram__T_3_data; // @[Decoupled.scala 209:16]
  wire [3:0] ram__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram__T_3_en; // @[Decoupled.scala 209:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 29:33]
  reg [3:0] deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  _T_1 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _T_5 = enq_ptr_value + 4'h1; // @[Counter.scala 39:22]
  wire  _GEN_9 = io_deq_ready ? 1'h0 : _T_1; // @[Decoupled.scala 240:27]
  wire  do_enq = empty ? _GEN_9 : _T_1; // @[Decoupled.scala 237:18]
  wire [3:0] _T_7 = deq_ptr_value + 4'h1; // @[Counter.scala 39:22]
  wire  do_deq = empty ? 1'h0 : _T_2; // @[Decoupled.scala 237:18]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  wire  _T_9 = ~empty; // @[Decoupled.scala 231:19]
  wire  _T_10 = ~full; // @[Decoupled.scala 232:19]
  assign ram__T_11_addr = deq_ptr_value;
  assign ram__T_11_data = ram[ram__T_11_addr]; // @[Decoupled.scala 209:16]
  assign ram__T_3_data = io_enq_bits;
  assign ram__T_3_addr = enq_ptr_value;
  assign ram__T_3_mask = 1'h1;
  assign ram__T_3_en = empty ? _GEN_9 : _T_1;
  assign io_enq_ready = io_deq_ready | _T_10; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = io_enq_valid | _T_9; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits = empty ? io_enq_bits : ram__T_11_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_3_en & ram__T_3_mask) begin
      ram[ram__T_3_addr] <= ram__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 4'h0;
    end else if (do_enq) begin
      enq_ptr_value <= _T_5;
    end
    if (reset) begin
      deq_ptr_value <= 4'h0;
    end else if (do_deq) begin
      deq_ptr_value <= _T_7;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _T_1;
        end
      end else begin
        maybe_full <= _T_1;
      end
    end
  end
endmodule
module memGenAccel(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_dataVals_field2_data,
  input  [63:0] io_in_bits_dataVals_field1_data,
  input  [63:0] io_in_bits_dataVals_field0_data,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_data_field1_data,
  output [31:0] io_events_bits_0,
  output [31:0] io_events_bits_1,
  output [31:0] io_events_bits_2,
  output [31:0] io_events_bits_3,
  output [31:0] io_events_bits_4,
  output [31:0] io_events_bits_5,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output        io_mem_b_ready,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [15:0] io_mem_ar_bits_len,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last
);
  wire  accel_clock; // @[memGenCacheShell.scala 24:22]
  wire  accel_reset; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_instruction_0_ready; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_instruction_0_valid; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_instruction_0_bits_addr; // @[memGenCacheShell.scala 24:22]
  wire [7:0] accel_io_instruction_0_bits_inst; // @[memGenCacheShell.scala 24:22]
  wire [63:0] accel_io_instruction_0_bits_data; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_resp_0_valid; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_resp_0_bits_addr; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_events_bits_0; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_events_bits_1; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_events_bits_2; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_events_bits_3; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_events_bits_4; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_events_bits_5; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_aw_ready; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_aw_valid; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_mem_aw_bits_addr; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_w_ready; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_w_valid; // @[memGenCacheShell.scala 24:22]
  wire [63:0] accel_io_mem_w_bits_data; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_b_ready; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_ar_ready; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_ar_valid; // @[memGenCacheShell.scala 24:22]
  wire [31:0] accel_io_mem_ar_bits_addr; // @[memGenCacheShell.scala 24:22]
  wire [15:0] accel_io_mem_ar_bits_len; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_r_ready; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_r_valid; // @[memGenCacheShell.scala 24:22]
  wire [63:0] accel_io_mem_r_bits_data; // @[memGenCacheShell.scala 24:22]
  wire  accel_io_mem_r_bits_last; // @[memGenCacheShell.scala 24:22]
  wire  outArb_io_in_0_ready; // @[memGenCacheShell.scala 33:22]
  wire  outArb_io_in_0_valid; // @[memGenCacheShell.scala 33:22]
  wire [31:0] outArb_io_in_0_bits; // @[memGenCacheShell.scala 33:22]
  wire  outArb_io_out_ready; // @[memGenCacheShell.scala 33:22]
  wire  outArb_io_out_valid; // @[memGenCacheShell.scala 33:22]
  wire [31:0] outArb_io_out_bits; // @[memGenCacheShell.scala 33:22]
  wire  outAddrQueue_0_clock; // @[memGenCacheShell.scala 36:19]
  wire  outAddrQueue_0_reset; // @[memGenCacheShell.scala 36:19]
  wire  outAddrQueue_0_io_enq_ready; // @[memGenCacheShell.scala 36:19]
  wire  outAddrQueue_0_io_enq_valid; // @[memGenCacheShell.scala 36:19]
  wire [31:0] outAddrQueue_0_io_enq_bits; // @[memGenCacheShell.scala 36:19]
  wire  outAddrQueue_0_io_deq_ready; // @[memGenCacheShell.scala 36:19]
  wire  outAddrQueue_0_io_deq_valid; // @[memGenCacheShell.scala 36:19]
  wire [31:0] outAddrQueue_0_io_deq_bits; // @[memGenCacheShell.scala 36:19]
  wire  _T = io_in_bits_dataVals_field0_data == 64'h4; // @[memGenCacheShell.scala 47:54]
  wire [63:0] _GEN_1 = _T ? 64'h0 : io_in_bits_dataVals_field0_data; // @[memGenCacheShell.scala 47:68]
  memGenTopLevel accel ( // @[memGenCacheShell.scala 24:22]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_instruction_0_ready(accel_io_instruction_0_ready),
    .io_instruction_0_valid(accel_io_instruction_0_valid),
    .io_instruction_0_bits_addr(accel_io_instruction_0_bits_addr),
    .io_instruction_0_bits_inst(accel_io_instruction_0_bits_inst),
    .io_instruction_0_bits_data(accel_io_instruction_0_bits_data),
    .io_resp_0_valid(accel_io_resp_0_valid),
    .io_resp_0_bits_addr(accel_io_resp_0_bits_addr),
    .io_events_bits_0(accel_io_events_bits_0),
    .io_events_bits_1(accel_io_events_bits_1),
    .io_events_bits_2(accel_io_events_bits_2),
    .io_events_bits_3(accel_io_events_bits_3),
    .io_events_bits_4(accel_io_events_bits_4),
    .io_events_bits_5(accel_io_events_bits_5),
    .io_mem_aw_ready(accel_io_mem_aw_ready),
    .io_mem_aw_valid(accel_io_mem_aw_valid),
    .io_mem_aw_bits_addr(accel_io_mem_aw_bits_addr),
    .io_mem_w_ready(accel_io_mem_w_ready),
    .io_mem_w_valid(accel_io_mem_w_valid),
    .io_mem_w_bits_data(accel_io_mem_w_bits_data),
    .io_mem_b_ready(accel_io_mem_b_ready),
    .io_mem_ar_ready(accel_io_mem_ar_ready),
    .io_mem_ar_valid(accel_io_mem_ar_valid),
    .io_mem_ar_bits_addr(accel_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(accel_io_mem_ar_bits_len),
    .io_mem_r_ready(accel_io_mem_r_ready),
    .io_mem_r_valid(accel_io_mem_r_valid),
    .io_mem_r_bits_data(accel_io_mem_r_bits_data),
    .io_mem_r_bits_last(accel_io_mem_r_bits_last)
  );
  Arbiter_6 outArb ( // @[memGenCacheShell.scala 33:22]
    .io_in_0_ready(outArb_io_in_0_ready),
    .io_in_0_valid(outArb_io_in_0_valid),
    .io_in_0_bits(outArb_io_in_0_bits),
    .io_out_ready(outArb_io_out_ready),
    .io_out_valid(outArb_io_out_valid),
    .io_out_bits(outArb_io_out_bits)
  );
  Queue_19 outAddrQueue_0 ( // @[memGenCacheShell.scala 36:19]
    .clock(outAddrQueue_0_clock),
    .reset(outAddrQueue_0_reset),
    .io_enq_ready(outAddrQueue_0_io_enq_ready),
    .io_enq_valid(outAddrQueue_0_io_enq_valid),
    .io_enq_bits(outAddrQueue_0_io_enq_bits),
    .io_deq_ready(outAddrQueue_0_io_deq_ready),
    .io_deq_valid(outAddrQueue_0_io_deq_valid),
    .io_deq_bits(outAddrQueue_0_io_deq_bits)
  );
  assign io_in_ready = accel_io_instruction_0_ready; // @[memGenCacheShell.scala 45:15 memGenCacheShell.scala 56:17]
  assign io_out_valid = outArb_io_out_valid; // @[memGenCacheShell.scala 74:16]
  assign io_out_bits_data_field1_data = outArb_io_out_bits; // @[memGenCacheShell.scala 75:35]
  assign io_events_bits_0 = accel_io_events_bits_0; // @[memGenCacheShell.scala 78:13]
  assign io_events_bits_1 = accel_io_events_bits_1; // @[memGenCacheShell.scala 78:13]
  assign io_events_bits_2 = accel_io_events_bits_2; // @[memGenCacheShell.scala 78:13]
  assign io_events_bits_3 = accel_io_events_bits_3; // @[memGenCacheShell.scala 78:13]
  assign io_events_bits_4 = accel_io_events_bits_4; // @[memGenCacheShell.scala 78:13]
  assign io_events_bits_5 = accel_io_events_bits_5; // @[memGenCacheShell.scala 78:13]
  assign io_mem_aw_valid = accel_io_mem_aw_valid; // @[memGenCacheShell.scala 80:10]
  assign io_mem_aw_bits_addr = accel_io_mem_aw_bits_addr; // @[memGenCacheShell.scala 80:10]
  assign io_mem_w_valid = accel_io_mem_w_valid; // @[memGenCacheShell.scala 80:10]
  assign io_mem_w_bits_data = accel_io_mem_w_bits_data; // @[memGenCacheShell.scala 80:10]
  assign io_mem_b_ready = accel_io_mem_b_ready; // @[memGenCacheShell.scala 80:10]
  assign io_mem_ar_valid = accel_io_mem_ar_valid; // @[memGenCacheShell.scala 80:10]
  assign io_mem_ar_bits_addr = accel_io_mem_ar_bits_addr; // @[memGenCacheShell.scala 80:10]
  assign io_mem_ar_bits_len = accel_io_mem_ar_bits_len; // @[memGenCacheShell.scala 80:10]
  assign io_mem_r_ready = accel_io_mem_r_ready; // @[memGenCacheShell.scala 80:10]
  assign accel_clock = clock;
  assign accel_reset = reset;
  assign accel_io_instruction_0_valid = io_in_valid; // @[memGenCacheShell.scala 39:41 memGenCacheShell.scala 57:41]
  assign accel_io_instruction_0_bits_addr = io_in_bits_dataVals_field1_data[31:0]; // @[memGenCacheShell.scala 41:45 memGenCacheShell.scala 58:45]
  assign accel_io_instruction_0_bits_inst = _GEN_1[7:0]; // @[memGenCacheShell.scala 40:45 memGenCacheShell.scala 50:47 memGenCacheShell.scala 52:49]
  assign accel_io_instruction_0_bits_data = io_in_bits_dataVals_field2_data; // @[memGenCacheShell.scala 42:45 memGenCacheShell.scala 59:45]
  assign accel_io_mem_aw_ready = io_mem_aw_ready; // @[memGenCacheShell.scala 80:10]
  assign accel_io_mem_w_ready = io_mem_w_ready; // @[memGenCacheShell.scala 80:10]
  assign accel_io_mem_ar_ready = io_mem_ar_ready; // @[memGenCacheShell.scala 80:10]
  assign accel_io_mem_r_valid = io_mem_r_valid; // @[memGenCacheShell.scala 80:10]
  assign accel_io_mem_r_bits_data = io_mem_r_bits_data; // @[memGenCacheShell.scala 80:10]
  assign accel_io_mem_r_bits_last = io_mem_r_bits_last; // @[memGenCacheShell.scala 80:10]
  assign outArb_io_in_0_valid = outAddrQueue_0_io_deq_valid; // @[memGenCacheShell.scala 71:21]
  assign outArb_io_in_0_bits = outAddrQueue_0_io_deq_bits; // @[memGenCacheShell.scala 71:21]
  assign outArb_io_out_ready = io_out_ready; // @[memGenCacheShell.scala 76:23]
  assign outAddrQueue_0_clock = clock;
  assign outAddrQueue_0_reset = reset;
  assign outAddrQueue_0_io_enq_valid = accel_io_resp_0_valid; // @[memGenCacheShell.scala 68:34]
  assign outAddrQueue_0_io_enq_bits = accel_io_resp_0_valid ? accel_io_resp_0_bits_addr : 32'h0; // @[memGenCacheShell.scala 67:33]
  assign outAddrQueue_0_io_deq_ready = outArb_io_in_0_ready; // @[memGenCacheShell.scala 71:21]
endmodule
module Queue_20(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_data
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_data [0:999999]; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_11_data; // @[Decoupled.scala 209:16]
  wire [19:0] ram_data__T_11_addr; // @[Decoupled.scala 209:16]
  wire [63:0] ram_data__T_3_data; // @[Decoupled.scala 209:16]
  wire [19:0] ram_data__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram_data__T_3_en; // @[Decoupled.scala 209:16]
  reg [19:0] enq_ptr_value; // @[Counter.scala 29:33]
  reg [19:0] deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  _T_1 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = enq_ptr_value == 20'hf423f; // @[Counter.scala 38:24]
  wire [19:0] _T_5 = enq_ptr_value + 20'h1; // @[Counter.scala 39:22]
  wire  _GEN_13 = io_deq_ready ? 1'h0 : _T_1; // @[Decoupled.scala 240:27]
  wire  do_enq = empty ? _GEN_13 : _T_1; // @[Decoupled.scala 237:18]
  wire  wrap_1 = deq_ptr_value == 20'hf423f; // @[Counter.scala 38:24]
  wire [19:0] _T_7 = deq_ptr_value + 20'h1; // @[Counter.scala 39:22]
  wire  do_deq = empty ? 1'h0 : _T_2; // @[Decoupled.scala 237:18]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  wire  _T_9 = ~empty; // @[Decoupled.scala 231:19]
  wire  _T_10 = ~full; // @[Decoupled.scala 232:19]
  assign ram_data__T_11_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_data__T_11_data = ram_data[ram_data__T_11_addr]; // @[Decoupled.scala 209:16]
  `else
  assign ram_data__T_11_data = ram_data__T_11_addr >= 20'hf4240 ? _RAND_1[63:0] : ram_data[ram_data__T_11_addr]; // @[Decoupled.scala 209:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_data__T_3_data = io_enq_bits_data;
  assign ram_data__T_3_addr = enq_ptr_value;
  assign ram_data__T_3_mask = 1'h1;
  assign ram_data__T_3_en = empty ? _GEN_13 : _T_1;
  assign io_enq_ready = io_deq_ready | _T_10; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = io_enq_valid | _T_9; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data__T_11_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {2{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1000000; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[19:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_data__T_3_en & ram_data__T_3_mask) begin
      ram_data[ram_data__T_3_addr] <= ram_data__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 20'h0;
    end else if (do_enq) begin
      if (wrap) begin
        enq_ptr_value <= 20'h0;
      end else begin
        enq_ptr_value <= _T_5;
      end
    end
    if (reset) begin
      deq_ptr_value <= 20'h0;
    end else if (do_deq) begin
      if (wrap_1) begin
        deq_ptr_value <= 20'h0;
      end else begin
        deq_ptr_value <= _T_7;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _T_1;
        end
      end else begin
        maybe_full <= _T_1;
      end
    end
  end
endmodule
module memGenDCRCacheShell(
  input         clock,
  input         reset,
  output        io_host_aw_ready,
  input         io_host_aw_valid,
  input  [31:0] io_host_aw_bits_addr,
  output        io_host_w_ready,
  input         io_host_w_valid,
  input  [63:0] io_host_w_bits_data,
  input         io_host_b_ready,
  output        io_host_b_valid,
  output        io_host_ar_ready,
  input         io_host_ar_valid,
  input  [31:0] io_host_ar_bits_addr,
  input         io_host_r_ready,
  output        io_host_r_valid,
  output [63:0] io_host_r_bits_data,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  output [31:0] io_mem_aw_bits_len,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output        io_mem_w_bits_last,
  output        io_mem_b_ready,
  input         io_mem_b_valid,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [31:0] io_mem_ar_bits_len,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  vcr_clock; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_reset; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_aw_ready; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_aw_valid; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_host_aw_bits_addr; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_w_ready; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_w_valid; // @[memGenDCRCacheShell.scala 37:19]
  wire [63:0] vcr_io_host_w_bits_data; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_b_ready; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_b_valid; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_ar_ready; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_ar_valid; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_host_ar_bits_addr; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_r_ready; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_host_r_valid; // @[memGenDCRCacheShell.scala 37:19]
  wire [63:0] vcr_io_host_r_bits_data; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_dcr_launch; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_dcr_finish; // @[memGenDCRCacheShell.scala 37:19]
  wire  vcr_io_dcr_ecnt_0_valid; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_0_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_1_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_2_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_3_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_4_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_5_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ecnt_6_bits; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_vals_0; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ptrs_1; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ptrs_2; // @[memGenDCRCacheShell.scala 37:19]
  wire [31:0] vcr_io_dcr_ptrs_3; // @[memGenDCRCacheShell.scala 37:19]
  wire  dmem_clock; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_reset; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_aw_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_aw_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_w_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_w_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_w_bits_last; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_b_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_b_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_ar_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_ar_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [31:0] dmem_io_mem_ar_bits_addr; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_r_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_r_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [63:0] dmem_io_mem_r_bits_data; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_mem_r_bits_last; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_0_cmd_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [31:0] dmem_io_dme_rd_0_cmd_bits_addr; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_0_data_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_0_data_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [63:0] dmem_io_dme_rd_0_data_bits; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_1_cmd_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [31:0] dmem_io_dme_rd_1_cmd_bits_addr; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_1_data_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_1_data_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [63:0] dmem_io_dme_rd_1_data_bits; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_2_cmd_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [31:0] dmem_io_dme_rd_2_cmd_bits_addr; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_2_data_ready; // @[memGenDCRCacheShell.scala 38:20]
  wire  dmem_io_dme_rd_2_data_valid; // @[memGenDCRCacheShell.scala 38:20]
  wire [63:0] dmem_io_dme_rd_2_data_bits; // @[memGenDCRCacheShell.scala 38:20]
  wire  accel_clock; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_reset; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_in_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_in_valid; // @[memGenDCRCacheShell.scala 40:21]
  wire [63:0] accel_io_in_bits_dataVals_field2_data; // @[memGenDCRCacheShell.scala 40:21]
  wire [63:0] accel_io_in_bits_dataVals_field1_data; // @[memGenDCRCacheShell.scala 40:21]
  wire [63:0] accel_io_in_bits_dataVals_field0_data; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_out_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_out_valid; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_out_bits_data_field1_data; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_events_bits_0; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_events_bits_1; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_events_bits_2; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_events_bits_3; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_events_bits_4; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_events_bits_5; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_aw_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_aw_valid; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_mem_aw_bits_addr; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_w_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_w_valid; // @[memGenDCRCacheShell.scala 40:21]
  wire [63:0] accel_io_mem_w_bits_data; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_b_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_ar_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_ar_valid; // @[memGenDCRCacheShell.scala 40:21]
  wire [31:0] accel_io_mem_ar_bits_addr; // @[memGenDCRCacheShell.scala 40:21]
  wire [15:0] accel_io_mem_ar_bits_len; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_r_ready; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_r_valid; // @[memGenDCRCacheShell.scala 40:21]
  wire [63:0] accel_io_mem_r_bits_data; // @[memGenDCRCacheShell.scala 40:21]
  wire  accel_io_mem_r_bits_last; // @[memGenDCRCacheShell.scala 40:21]
  wire  inputQ_0_clock; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_0_reset; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_0_io_enq_ready; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_0_io_enq_valid; // @[memGenDCRCacheShell.scala 113:25]
  wire [63:0] inputQ_0_io_enq_bits_data; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_0_io_deq_ready; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_0_io_deq_valid; // @[memGenDCRCacheShell.scala 113:25]
  wire [63:0] inputQ_0_io_deq_bits_data; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_1_clock; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_1_reset; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_1_io_enq_ready; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_1_io_enq_valid; // @[memGenDCRCacheShell.scala 113:25]
  wire [63:0] inputQ_1_io_enq_bits_data; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_1_io_deq_ready; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_1_io_deq_valid; // @[memGenDCRCacheShell.scala 113:25]
  wire [63:0] inputQ_1_io_deq_bits_data; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_2_clock; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_2_reset; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_2_io_enq_ready; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_2_io_enq_valid; // @[memGenDCRCacheShell.scala 113:25]
  wire [63:0] inputQ_2_io_enq_bits_data; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_2_io_deq_ready; // @[memGenDCRCacheShell.scala 113:25]
  wire  inputQ_2_io_deq_valid; // @[memGenDCRCacheShell.scala 113:25]
  wire [63:0] inputQ_2_io_deq_bits_data; // @[memGenDCRCacheShell.scala 113:25]
  reg [2:0] state; // @[memGenDCRCacheShell.scala 46:22]
  reg [31:0] cycles; // @[memGenDCRCacheShell.scala 47:23]
  wire  last = state == 3'h5; // @[memGenDCRCacheShell.scala 48:20]
  wire  is_busy = state == 3'h2; // @[memGenDCRCacheShell.scala 49:23]
  reg [31:0] lastCycle; // @[memGenDCRCacheShell.scala 53:21]
  reg [14:0] cycle; // @[Counter.scala 29:33]
  wire  _T_1 = cycle == 15'h752f; // @[Counter.scala 38:24]
  wire [14:0] _T_3 = cycle + 15'h1; // @[Counter.scala 39:22]
  wire  stopSim = last & _T_1; // @[Counter.scala 67:17]
  wire  _T_4 = state == 3'h0; // @[memGenDCRCacheShell.scala 74:128]
  reg [63:0] vals_0; // @[Reg.scala 27:20]
  wire  _T_75 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_76 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_77 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_78 = ~inputQ_0_io_deq_valid; // @[memGenDCRCacheShell.scala 169:37]
  wire  _T_79 = inputQ_0_io_deq_bits_data == 64'h2; // @[memGenDCRCacheShell.scala 171:54]
  wire  _T_82 = inputQ_0_io_deq_bits_data == 64'h4; // @[memGenDCRCacheShell.scala 174:53]
  wire  _T_83 = accel_io_in_ready & accel_io_in_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_28 = _T_82 | _T_83; // @[memGenDCRCacheShell.scala 174:66]
  wire  _GEN_31 = _T_79 ? 1'h0 : _GEN_28; // @[memGenDCRCacheShell.scala 171:68]
  wire  _GEN_34 = _T_78 ? 1'h0 : _GEN_31; // @[memGenDCRCacheShell.scala 169:93]
  wire  _T_86 = 3'h4 == state; // @[Conditional.scala 37:30]
  reg [19:0] ackCounter; // @[Counter.scala 29:33]
  wire [63:0] _GEN_112 = {{44'd0}, ackCounter}; // @[memGenDCRCacheShell.scala 186:26]
  wire  _T_87 = _GEN_112 >= inputQ_2_io_deq_bits_data; // @[memGenDCRCacheShell.scala 186:26]
  wire  _GEN_41 = _T_86 & _T_87; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_77 ? _GEN_34 : _GEN_41; // @[Conditional.scala 39:67]
  wire  _GEN_47 = _T_76 ? 1'h0 : _GEN_43; // @[Conditional.scala 39:67]
  wire  _T_19 = ackCounter == 20'hf423f; // @[Counter.scala 38:24]
  wire [19:0] _T_21 = ackCounter + 20'h1; // @[Counter.scala 39:22]
  wire  _GEN_45 = _T_77 ? 1'h0 : _GEN_41; // @[Conditional.scala 39:67]
  wire  _GEN_49 = _T_76 ? 1'h0 : _GEN_45; // @[Conditional.scala 39:67]
  wire  resetAckCounter = _T_75 ? 1'h0 : _GEN_49; // @[Conditional.scala 40:58]
  reg [31:0] fillCounter; // @[memGenDCRCacheShell.scala 79:28]
  wire  _T_22 = dmem_io_mem_r_ready & dmem_io_mem_r_valid; // @[Decoupled.scala 40:37]
  reg [31:0] _T_29; // @[memGenDCRCacheShell.scala 92:22]
  wire [63:0] _T_30 = vals_0 / 64'h1; // @[memGenDCRCacheShell.scala 92:50]
  wire [63:0] _T_32 = _T_30 - 64'h1; // @[memGenDCRCacheShell.scala 92:61]
  wire [63:0] _GEN_113 = {{32'd0}, _T_29}; // @[memGenDCRCacheShell.scala 92:36]
  wire  fillWrap = _GEN_113 == _T_32; // @[memGenDCRCacheShell.scala 92:36]
  wire  _T_23 = fillWrap & _T_22; // @[memGenDCRCacheShell.scala 85:18]
  wire  _T_24 = _T_23 & dmem_io_mem_r_bits_last; // @[memGenDCRCacheShell.scala 85:42]
  wire  _T_26 = _T_22 & dmem_io_mem_r_bits_last; // @[memGenDCRCacheShell.scala 87:35]
  wire [31:0] _T_28 = fillCounter + 32'h1; // @[memGenDCRCacheShell.scala 88:32]
  reg [1:0] numQ; // @[Counter.scala 29:33]
  wire [1:0] _T_40 = numQ + 2'h1; // @[Counter.scala 39:22]
  wire  _T_43 = numQ == 2'h2; // @[memGenDCRCacheShell.scala 95:72]
  wire  _T_44 = _T_26 & _T_43; // @[memGenDCRCacheShell.scala 95:64]
  wire  goToBusy = _T_44 & fillWrap; // @[memGenDCRCacheShell.scala 95:80]
  wire [31:0] _T_47 = cycles + 32'h1; // @[memGenDCRCacheShell.scala 100:22]
  wire  _T_48 = accel_io_out_ready & accel_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_50 = ~reset; // @[memGenDCRCacheShell.scala 107:13]
  wire [32:0] _T_53 = fillCounter * 32'h1; // @[memGenDCRCacheShell.scala 120:79]
  wire [36:0] _T_54 = _T_53 * 33'h8; // @[memGenDCRCacheShell.scala 120:89]
  wire [36:0] _GEN_114 = {{5'd0}, vcr_io_dcr_ptrs_1}; // @[memGenDCRCacheShell.scala 120:65]
  wire [36:0] _T_56 = _GEN_114 + _T_54; // @[memGenDCRCacheShell.scala 120:65]
  wire [36:0] _GEN_115 = {{5'd0}, vcr_io_dcr_ptrs_2}; // @[memGenDCRCacheShell.scala 120:65]
  wire [36:0] _T_61 = _GEN_115 + _T_54; // @[memGenDCRCacheShell.scala 120:65]
  wire [36:0] _GEN_116 = {{5'd0}, vcr_io_dcr_ptrs_3}; // @[memGenDCRCacheShell.scala 120:65]
  wire [36:0] _T_66 = _GEN_116 + _T_54; // @[memGenDCRCacheShell.scala 120:65]
  wire  _T_68 = state == 3'h1; // @[memGenDCRCacheShell.scala 131:47]
  wire  _GEN_117 = 2'h0 == numQ; // @[memGenDCRCacheShell.scala 131:36]
  wire  _GEN_118 = 2'h1 == numQ; // @[memGenDCRCacheShell.scala 131:36]
  wire  _GEN_119 = 2'h2 == numQ; // @[memGenDCRCacheShell.scala 131:36]
  wire  _T_72 = is_busy | last; // @[memGenDCRCacheShell.scala 151:33]
  wire  _T_73 = state == 3'h4; // @[memGenDCRCacheShell.scala 151:59]
  wire  _GEN_29 = _T_82 ? 1'h0 : 1'h1; // @[memGenDCRCacheShell.scala 174:66]
  wire  _GEN_32 = _T_79 ? 1'h0 : _GEN_29; // @[memGenDCRCacheShell.scala 171:68]
  wire  _GEN_35 = _T_78 ? 1'h0 : _GEN_32; // @[memGenDCRCacheShell.scala 169:93]
  wire  _T_88 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_44 = _T_77 & _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_48 = _T_76 ? 1'h0 : _GEN_44; // @[Conditional.scala 39:67]
  wire  _GEN_123 = ~_T_75; // @[memGenDCRCacheShell.scala 173:17]
  wire  _GEN_124 = ~_T_76; // @[memGenDCRCacheShell.scala 173:17]
  wire  _GEN_125 = _GEN_123 & _GEN_124; // @[memGenDCRCacheShell.scala 173:17]
  wire  _GEN_126 = _GEN_125 & _T_77; // @[memGenDCRCacheShell.scala 173:17]
  wire  _GEN_127 = ~_T_78; // @[memGenDCRCacheShell.scala 173:17]
  wire  _GEN_128 = _GEN_126 & _GEN_127; // @[memGenDCRCacheShell.scala 173:17]
  wire  _GEN_129 = _GEN_128 & _T_79; // @[memGenDCRCacheShell.scala 173:17]
  wire  _GEN_136 = ~_T_79; // @[memGenDCRCacheShell.scala 179:21]
  wire  _GEN_137 = _GEN_128 & _GEN_136; // @[memGenDCRCacheShell.scala 179:21]
  wire  _GEN_138 = ~_T_82; // @[memGenDCRCacheShell.scala 179:21]
  wire  _GEN_139 = _GEN_137 & _GEN_138; // @[memGenDCRCacheShell.scala 179:21]
  wire  _GEN_140 = _GEN_139 & _T_83; // @[memGenDCRCacheShell.scala 179:21]
  DCR vcr ( // @[memGenDCRCacheShell.scala 37:19]
    .clock(vcr_clock),
    .reset(vcr_reset),
    .io_host_aw_ready(vcr_io_host_aw_ready),
    .io_host_aw_valid(vcr_io_host_aw_valid),
    .io_host_aw_bits_addr(vcr_io_host_aw_bits_addr),
    .io_host_w_ready(vcr_io_host_w_ready),
    .io_host_w_valid(vcr_io_host_w_valid),
    .io_host_w_bits_data(vcr_io_host_w_bits_data),
    .io_host_b_ready(vcr_io_host_b_ready),
    .io_host_b_valid(vcr_io_host_b_valid),
    .io_host_ar_ready(vcr_io_host_ar_ready),
    .io_host_ar_valid(vcr_io_host_ar_valid),
    .io_host_ar_bits_addr(vcr_io_host_ar_bits_addr),
    .io_host_r_ready(vcr_io_host_r_ready),
    .io_host_r_valid(vcr_io_host_r_valid),
    .io_host_r_bits_data(vcr_io_host_r_bits_data),
    .io_dcr_launch(vcr_io_dcr_launch),
    .io_dcr_finish(vcr_io_dcr_finish),
    .io_dcr_ecnt_0_valid(vcr_io_dcr_ecnt_0_valid),
    .io_dcr_ecnt_0_bits(vcr_io_dcr_ecnt_0_bits),
    .io_dcr_ecnt_1_bits(vcr_io_dcr_ecnt_1_bits),
    .io_dcr_ecnt_2_bits(vcr_io_dcr_ecnt_2_bits),
    .io_dcr_ecnt_3_bits(vcr_io_dcr_ecnt_3_bits),
    .io_dcr_ecnt_4_bits(vcr_io_dcr_ecnt_4_bits),
    .io_dcr_ecnt_5_bits(vcr_io_dcr_ecnt_5_bits),
    .io_dcr_ecnt_6_bits(vcr_io_dcr_ecnt_6_bits),
    .io_dcr_vals_0(vcr_io_dcr_vals_0),
    .io_dcr_ptrs_1(vcr_io_dcr_ptrs_1),
    .io_dcr_ptrs_2(vcr_io_dcr_ptrs_2),
    .io_dcr_ptrs_3(vcr_io_dcr_ptrs_3)
  );
  DME dmem ( // @[memGenDCRCacheShell.scala 38:20]
    .clock(dmem_clock),
    .reset(dmem_reset),
    .io_mem_aw_ready(dmem_io_mem_aw_ready),
    .io_mem_aw_valid(dmem_io_mem_aw_valid),
    .io_mem_w_ready(dmem_io_mem_w_ready),
    .io_mem_w_valid(dmem_io_mem_w_valid),
    .io_mem_w_bits_last(dmem_io_mem_w_bits_last),
    .io_mem_b_ready(dmem_io_mem_b_ready),
    .io_mem_b_valid(dmem_io_mem_b_valid),
    .io_mem_ar_ready(dmem_io_mem_ar_ready),
    .io_mem_ar_valid(dmem_io_mem_ar_valid),
    .io_mem_ar_bits_addr(dmem_io_mem_ar_bits_addr),
    .io_mem_r_ready(dmem_io_mem_r_ready),
    .io_mem_r_valid(dmem_io_mem_r_valid),
    .io_mem_r_bits_data(dmem_io_mem_r_bits_data),
    .io_mem_r_bits_last(dmem_io_mem_r_bits_last),
    .io_dme_rd_0_cmd_valid(dmem_io_dme_rd_0_cmd_valid),
    .io_dme_rd_0_cmd_bits_addr(dmem_io_dme_rd_0_cmd_bits_addr),
    .io_dme_rd_0_data_ready(dmem_io_dme_rd_0_data_ready),
    .io_dme_rd_0_data_valid(dmem_io_dme_rd_0_data_valid),
    .io_dme_rd_0_data_bits(dmem_io_dme_rd_0_data_bits),
    .io_dme_rd_1_cmd_valid(dmem_io_dme_rd_1_cmd_valid),
    .io_dme_rd_1_cmd_bits_addr(dmem_io_dme_rd_1_cmd_bits_addr),
    .io_dme_rd_1_data_ready(dmem_io_dme_rd_1_data_ready),
    .io_dme_rd_1_data_valid(dmem_io_dme_rd_1_data_valid),
    .io_dme_rd_1_data_bits(dmem_io_dme_rd_1_data_bits),
    .io_dme_rd_2_cmd_valid(dmem_io_dme_rd_2_cmd_valid),
    .io_dme_rd_2_cmd_bits_addr(dmem_io_dme_rd_2_cmd_bits_addr),
    .io_dme_rd_2_data_ready(dmem_io_dme_rd_2_data_ready),
    .io_dme_rd_2_data_valid(dmem_io_dme_rd_2_data_valid),
    .io_dme_rd_2_data_bits(dmem_io_dme_rd_2_data_bits)
  );
  memGenAccel accel ( // @[memGenDCRCacheShell.scala 40:21]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_in_ready(accel_io_in_ready),
    .io_in_valid(accel_io_in_valid),
    .io_in_bits_dataVals_field2_data(accel_io_in_bits_dataVals_field2_data),
    .io_in_bits_dataVals_field1_data(accel_io_in_bits_dataVals_field1_data),
    .io_in_bits_dataVals_field0_data(accel_io_in_bits_dataVals_field0_data),
    .io_out_ready(accel_io_out_ready),
    .io_out_valid(accel_io_out_valid),
    .io_out_bits_data_field1_data(accel_io_out_bits_data_field1_data),
    .io_events_bits_0(accel_io_events_bits_0),
    .io_events_bits_1(accel_io_events_bits_1),
    .io_events_bits_2(accel_io_events_bits_2),
    .io_events_bits_3(accel_io_events_bits_3),
    .io_events_bits_4(accel_io_events_bits_4),
    .io_events_bits_5(accel_io_events_bits_5),
    .io_mem_aw_ready(accel_io_mem_aw_ready),
    .io_mem_aw_valid(accel_io_mem_aw_valid),
    .io_mem_aw_bits_addr(accel_io_mem_aw_bits_addr),
    .io_mem_w_ready(accel_io_mem_w_ready),
    .io_mem_w_valid(accel_io_mem_w_valid),
    .io_mem_w_bits_data(accel_io_mem_w_bits_data),
    .io_mem_b_ready(accel_io_mem_b_ready),
    .io_mem_ar_ready(accel_io_mem_ar_ready),
    .io_mem_ar_valid(accel_io_mem_ar_valid),
    .io_mem_ar_bits_addr(accel_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(accel_io_mem_ar_bits_len),
    .io_mem_r_ready(accel_io_mem_r_ready),
    .io_mem_r_valid(accel_io_mem_r_valid),
    .io_mem_r_bits_data(accel_io_mem_r_bits_data),
    .io_mem_r_bits_last(accel_io_mem_r_bits_last)
  );
  Queue_20 inputQ_0 ( // @[memGenDCRCacheShell.scala 113:25]
    .clock(inputQ_0_clock),
    .reset(inputQ_0_reset),
    .io_enq_ready(inputQ_0_io_enq_ready),
    .io_enq_valid(inputQ_0_io_enq_valid),
    .io_enq_bits_data(inputQ_0_io_enq_bits_data),
    .io_deq_ready(inputQ_0_io_deq_ready),
    .io_deq_valid(inputQ_0_io_deq_valid),
    .io_deq_bits_data(inputQ_0_io_deq_bits_data)
  );
  Queue_20 inputQ_1 ( // @[memGenDCRCacheShell.scala 113:25]
    .clock(inputQ_1_clock),
    .reset(inputQ_1_reset),
    .io_enq_ready(inputQ_1_io_enq_ready),
    .io_enq_valid(inputQ_1_io_enq_valid),
    .io_enq_bits_data(inputQ_1_io_enq_bits_data),
    .io_deq_ready(inputQ_1_io_deq_ready),
    .io_deq_valid(inputQ_1_io_deq_valid),
    .io_deq_bits_data(inputQ_1_io_deq_bits_data)
  );
  Queue_20 inputQ_2 ( // @[memGenDCRCacheShell.scala 113:25]
    .clock(inputQ_2_clock),
    .reset(inputQ_2_reset),
    .io_enq_ready(inputQ_2_io_enq_ready),
    .io_enq_valid(inputQ_2_io_enq_valid),
    .io_enq_bits_data(inputQ_2_io_enq_bits_data),
    .io_deq_ready(inputQ_2_io_deq_ready),
    .io_deq_valid(inputQ_2_io_deq_valid),
    .io_deq_bits_data(inputQ_2_io_deq_bits_data)
  );
  assign io_host_aw_ready = vcr_io_host_aw_ready; // @[memGenDCRCacheShell.scala 210:11]
  assign io_host_w_ready = vcr_io_host_w_ready; // @[memGenDCRCacheShell.scala 210:11]
  assign io_host_b_valid = vcr_io_host_b_valid; // @[memGenDCRCacheShell.scala 210:11]
  assign io_host_ar_ready = vcr_io_host_ar_ready; // @[memGenDCRCacheShell.scala 210:11]
  assign io_host_r_valid = vcr_io_host_r_valid; // @[memGenDCRCacheShell.scala 210:11]
  assign io_host_r_bits_data = vcr_io_host_r_bits_data; // @[memGenDCRCacheShell.scala 210:11]
  assign io_mem_aw_valid = _T_68 ? dmem_io_mem_aw_valid : accel_io_mem_aw_valid; // @[memGenDCRCacheShell.scala 203:12 memGenDCRCacheShell.scala 206:13]
  assign io_mem_aw_bits_addr = _T_68 ? 32'h0 : accel_io_mem_aw_bits_addr; // @[memGenDCRCacheShell.scala 203:12 memGenDCRCacheShell.scala 206:13]
  assign io_mem_aw_bits_len = _T_68 ? 32'h0 : 32'h1; // @[memGenDCRCacheShell.scala 203:12 memGenDCRCacheShell.scala 206:13]
  assign io_mem_w_valid = _T_68 ? 1'h0 : accel_io_mem_w_valid; // @[memGenDCRCacheShell.scala 203:12 memGenDCRCacheShell.scala 206:13]
  assign io_mem_w_bits_data = _T_68 ? 64'h0 : accel_io_mem_w_bits_data; // @[memGenDCRCacheShell.scala 203:12 memGenDCRCacheShell.scala 206:13]
  assign io_mem_w_bits_last = _T_68 & dmem_io_mem_w_bits_last; // @[memGenDCRCacheShell.scala 203:12 memGenDCRCacheShell.scala 206:13]
  assign io_mem_b_ready = _T_68 ? dmem_io_mem_b_ready : accel_io_mem_b_ready; // @[memGenDCRCacheShell.scala 203:12 memGenDCRCacheShell.scala 206:13]
  assign io_mem_ar_valid = _T_68 ? dmem_io_mem_ar_valid : accel_io_mem_ar_valid; // @[memGenDCRCacheShell.scala 203:12 memGenDCRCacheShell.scala 206:13]
  assign io_mem_ar_bits_addr = _T_68 ? dmem_io_mem_ar_bits_addr : accel_io_mem_ar_bits_addr; // @[memGenDCRCacheShell.scala 203:12 memGenDCRCacheShell.scala 206:13]
  assign io_mem_ar_bits_len = _T_68 ? 32'h0 : {{16'd0}, accel_io_mem_ar_bits_len}; // @[memGenDCRCacheShell.scala 203:12 memGenDCRCacheShell.scala 206:13]
  assign io_mem_r_ready = _T_68 ? dmem_io_mem_r_ready : accel_io_mem_r_ready; // @[memGenDCRCacheShell.scala 203:12 memGenDCRCacheShell.scala 206:13]
  assign vcr_clock = clock;
  assign vcr_reset = reset;
  assign vcr_io_host_aw_valid = io_host_aw_valid; // @[memGenDCRCacheShell.scala 210:11]
  assign vcr_io_host_aw_bits_addr = io_host_aw_bits_addr; // @[memGenDCRCacheShell.scala 210:11]
  assign vcr_io_host_w_valid = io_host_w_valid; // @[memGenDCRCacheShell.scala 210:11]
  assign vcr_io_host_w_bits_data = io_host_w_bits_data; // @[memGenDCRCacheShell.scala 210:11]
  assign vcr_io_host_b_ready = io_host_b_ready; // @[memGenDCRCacheShell.scala 210:11]
  assign vcr_io_host_ar_valid = io_host_ar_valid; // @[memGenDCRCacheShell.scala 210:11]
  assign vcr_io_host_ar_bits_addr = io_host_ar_bits_addr; // @[memGenDCRCacheShell.scala 210:11]
  assign vcr_io_host_r_ready = io_host_r_ready; // @[memGenDCRCacheShell.scala 210:11]
  assign vcr_io_dcr_finish = last & stopSim; // @[memGenDCRCacheShell.scala 200:21]
  assign vcr_io_dcr_ecnt_0_valid = state == 3'h5; // @[memGenDCRCacheShell.scala 103:27]
  assign vcr_io_dcr_ecnt_0_bits = lastCycle; // @[memGenDCRCacheShell.scala 104:26]
  assign vcr_io_dcr_ecnt_1_bits = accel_io_events_bits_0; // @[memGenDCRCacheShell.scala 63:31]
  assign vcr_io_dcr_ecnt_2_bits = accel_io_events_bits_1; // @[memGenDCRCacheShell.scala 63:31]
  assign vcr_io_dcr_ecnt_3_bits = accel_io_events_bits_2; // @[memGenDCRCacheShell.scala 63:31]
  assign vcr_io_dcr_ecnt_4_bits = accel_io_events_bits_3; // @[memGenDCRCacheShell.scala 63:31]
  assign vcr_io_dcr_ecnt_5_bits = accel_io_events_bits_4; // @[memGenDCRCacheShell.scala 63:31]
  assign vcr_io_dcr_ecnt_6_bits = accel_io_events_bits_5; // @[memGenDCRCacheShell.scala 63:31]
  assign dmem_clock = clock;
  assign dmem_reset = reset;
  assign dmem_io_mem_aw_ready = io_mem_aw_ready; // @[memGenDCRCacheShell.scala 203:12]
  assign dmem_io_mem_w_ready = io_mem_w_ready; // @[memGenDCRCacheShell.scala 203:12]
  assign dmem_io_mem_b_valid = io_mem_b_valid; // @[memGenDCRCacheShell.scala 203:12]
  assign dmem_io_mem_ar_ready = io_mem_ar_ready; // @[memGenDCRCacheShell.scala 203:12]
  assign dmem_io_mem_r_valid = io_mem_r_valid; // @[memGenDCRCacheShell.scala 203:12]
  assign dmem_io_mem_r_bits_data = io_mem_r_bits_data; // @[memGenDCRCacheShell.scala 203:12]
  assign dmem_io_mem_r_bits_last = io_mem_r_bits_last; // @[memGenDCRCacheShell.scala 203:12]
  assign dmem_io_dme_rd_0_cmd_valid = _GEN_117 & _T_68; // @[memGenDCRCacheShell.scala 122:39 memGenDCRCacheShell.scala 131:36]
  assign dmem_io_dme_rd_0_cmd_bits_addr = _T_56[31:0]; // @[memGenDCRCacheShell.scala 120:39]
  assign dmem_io_dme_rd_0_data_ready = inputQ_0_io_enq_ready; // @[memGenDCRCacheShell.scala 123:36]
  assign dmem_io_dme_rd_1_cmd_valid = _GEN_118 & _T_68; // @[memGenDCRCacheShell.scala 122:39 memGenDCRCacheShell.scala 131:36]
  assign dmem_io_dme_rd_1_cmd_bits_addr = _T_61[31:0]; // @[memGenDCRCacheShell.scala 120:39]
  assign dmem_io_dme_rd_1_data_ready = inputQ_1_io_enq_ready; // @[memGenDCRCacheShell.scala 123:36]
  assign dmem_io_dme_rd_2_cmd_valid = _GEN_119 & _T_68; // @[memGenDCRCacheShell.scala 122:39 memGenDCRCacheShell.scala 131:36]
  assign dmem_io_dme_rd_2_cmd_bits_addr = _T_66[31:0]; // @[memGenDCRCacheShell.scala 120:39]
  assign dmem_io_dme_rd_2_data_ready = inputQ_2_io_enq_ready; // @[memGenDCRCacheShell.scala 123:36]
  assign accel_clock = clock;
  assign accel_reset = reset;
  assign accel_io_in_valid = _T_75 ? 1'h0 : _GEN_48; // @[memGenDCRCacheShell.scala 150:21 memGenDCRCacheShell.scala 177:31]
  assign accel_io_in_bits_dataVals_field2_data = inputQ_2_io_deq_bits_data; // @[memGenDCRCacheShell.scala 144:47 memGenDCRCacheShell.scala 146:42]
  assign accel_io_in_bits_dataVals_field1_data = inputQ_1_io_deq_bits_data; // @[memGenDCRCacheShell.scala 140:45]
  assign accel_io_in_bits_dataVals_field0_data = inputQ_0_io_deq_bits_data; // @[memGenDCRCacheShell.scala 140:45]
  assign accel_io_out_ready = _T_72 | _T_73; // @[memGenDCRCacheShell.scala 151:22]
  assign accel_io_mem_aw_ready = io_mem_aw_ready; // @[memGenDCRCacheShell.scala 206:13]
  assign accel_io_mem_w_ready = io_mem_w_ready; // @[memGenDCRCacheShell.scala 206:13]
  assign accel_io_mem_ar_ready = io_mem_ar_ready; // @[memGenDCRCacheShell.scala 206:13]
  assign accel_io_mem_r_valid = io_mem_r_valid; // @[memGenDCRCacheShell.scala 206:13]
  assign accel_io_mem_r_bits_data = io_mem_r_bits_data; // @[memGenDCRCacheShell.scala 206:13]
  assign accel_io_mem_r_bits_last = io_mem_r_bits_last; // @[memGenDCRCacheShell.scala 206:13]
  assign inputQ_0_clock = clock;
  assign inputQ_0_reset = reset;
  assign inputQ_0_io_enq_valid = dmem_io_dme_rd_0_data_valid; // @[memGenDCRCacheShell.scala 126:30]
  assign inputQ_0_io_enq_bits_data = dmem_io_dme_rd_0_data_bits; // @[memGenDCRCacheShell.scala 125:29]
  assign inputQ_0_io_deq_ready = _T_75 ? 1'h0 : _GEN_47; // @[memGenDCRCacheShell.scala 127:30]
  assign inputQ_1_clock = clock;
  assign inputQ_1_reset = reset;
  assign inputQ_1_io_enq_valid = dmem_io_dme_rd_1_data_valid; // @[memGenDCRCacheShell.scala 126:30]
  assign inputQ_1_io_enq_bits_data = dmem_io_dme_rd_1_data_bits; // @[memGenDCRCacheShell.scala 125:29]
  assign inputQ_1_io_deq_ready = _T_75 ? 1'h0 : _GEN_47; // @[memGenDCRCacheShell.scala 127:30]
  assign inputQ_2_clock = clock;
  assign inputQ_2_reset = reset;
  assign inputQ_2_io_enq_valid = dmem_io_dme_rd_2_data_valid; // @[memGenDCRCacheShell.scala 126:30]
  assign inputQ_2_io_enq_bits_data = dmem_io_dme_rd_2_data_bits; // @[memGenDCRCacheShell.scala 125:29]
  assign inputQ_2_io_deq_ready = _T_75 ? 1'h0 : _GEN_47; // @[memGenDCRCacheShell.scala 127:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  cycles = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  lastCycle = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  cycle = _RAND_3[14:0];
  _RAND_4 = {2{`RANDOM}};
  vals_0 = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  ackCounter = _RAND_5[19:0];
  _RAND_6 = {1{`RANDOM}};
  fillCounter = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  _T_29 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  numQ = _RAND_8[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else if (_T_75) begin
      if (vcr_io_dcr_launch) begin
        state <= 3'h1;
      end
    end else if (_T_76) begin
      if (goToBusy) begin
        state <= 3'h2;
      end
    end else if (_T_77) begin
      if (_T_78) begin
        state <= 3'h5;
      end else if (_T_79) begin
        state <= 3'h4;
      end
    end else if (_T_86) begin
      if (_T_87) begin
        state <= 3'h2;
      end
    end else if (_T_88) begin
      if (stopSim) begin
        state <= 3'h0;
      end
    end
    if (reset) begin
      cycles <= 32'h0;
    end else if (goToBusy) begin
      cycles <= 32'h0;
    end else begin
      cycles <= _T_47;
    end
    if (_T_48) begin
      lastCycle <= cycles;
    end
    if (reset) begin
      cycle <= 15'h0;
    end else if (last) begin
      if (_T_1) begin
        cycle <= 15'h0;
      end else begin
        cycle <= _T_3;
      end
    end
    if (reset) begin
      vals_0 <= 64'h0;
    end else if (_T_4) begin
      vals_0 <= {{32'd0}, vcr_io_dcr_vals_0};
    end
    if (reset) begin
      ackCounter <= 20'h0;
    end else if (resetAckCounter) begin
      ackCounter <= 20'h0;
    end else if (accel_io_out_valid) begin
      if (_T_19) begin
        ackCounter <= 20'h0;
      end else begin
        ackCounter <= _T_21;
      end
    end
    if (reset) begin
      fillCounter <= 32'h0;
    end else if (_T_24) begin
      fillCounter <= 32'h0;
    end else if (_T_26) begin
      fillCounter <= _T_28;
    end
    _T_29 <= fillCounter;
    if (reset) begin
      numQ <= 2'h0;
    end else if (_T_24) begin
      numQ <= _T_40;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_48 & _T_50) begin
          $fwrite(32'h80000002,"Data back for addr %d cycle %d \n",accel_io_out_bits_data_field1_data,cycles); // @[memGenDCRCacheShell.scala 107:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_48 & _T_50) begin
          $fwrite(32'h80000002,"ackCounter :%d\n",ackCounter); // @[memGenDCRCacheShell.scala 108:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_129 & _T_50) begin
          $fwrite(32'h80000002,"Ack \n"); // @[memGenDCRCacheShell.scala 173:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_140 & _T_50) begin
          $fwrite(32'h80000002,"\nInst : %d for addr %d with data %d cycle %d \n",accel_io_in_bits_dataVals_field0_data,accel_io_in_bits_dataVals_field1_data,accel_io_in_bits_dataVals_field2_data,cycles); // @[memGenDCRCacheShell.scala 179:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module DandelionSimDCRAccel(
  input   clock,
  input   reset,
  input   sim_clock,
  output  sim_wait
);
  wire  sim_shell_clock; // @[DCRAccel.scala 52:25]
  wire  sim_shell_reset; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_aw_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_aw_valid; // @[DCRAccel.scala 52:25]
  wire [31:0] sim_shell_mem_aw_bits_addr; // @[DCRAccel.scala 52:25]
  wire [31:0] sim_shell_mem_aw_bits_len; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_w_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_w_valid; // @[DCRAccel.scala 52:25]
  wire [63:0] sim_shell_mem_w_bits_data; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_w_bits_last; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_b_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_b_valid; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_ar_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_ar_valid; // @[DCRAccel.scala 52:25]
  wire [31:0] sim_shell_mem_ar_bits_addr; // @[DCRAccel.scala 52:25]
  wire [31:0] sim_shell_mem_ar_bits_len; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_r_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_r_valid; // @[DCRAccel.scala 52:25]
  wire [63:0] sim_shell_mem_r_bits_data; // @[DCRAccel.scala 52:25]
  wire  sim_shell_mem_r_bits_last; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_aw_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_aw_valid; // @[DCRAccel.scala 52:25]
  wire [31:0] sim_shell_host_aw_bits_addr; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_w_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_w_valid; // @[DCRAccel.scala 52:25]
  wire [63:0] sim_shell_host_w_bits_data; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_b_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_b_valid; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_ar_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_ar_valid; // @[DCRAccel.scala 52:25]
  wire [31:0] sim_shell_host_ar_bits_addr; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_r_ready; // @[DCRAccel.scala 52:25]
  wire  sim_shell_host_r_valid; // @[DCRAccel.scala 52:25]
  wire [63:0] sim_shell_host_r_bits_data; // @[DCRAccel.scala 52:25]
  wire  sim_shell_sim_clock; // @[DCRAccel.scala 52:25]
  wire  sim_shell_sim_wait; // @[DCRAccel.scala 52:25]
  wire  shell_clock; // @[DCRAccel.scala 53:21]
  wire  shell_reset; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_aw_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_aw_valid; // @[DCRAccel.scala 53:21]
  wire [31:0] shell_io_host_aw_bits_addr; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_w_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_w_valid; // @[DCRAccel.scala 53:21]
  wire [63:0] shell_io_host_w_bits_data; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_b_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_b_valid; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_ar_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_ar_valid; // @[DCRAccel.scala 53:21]
  wire [31:0] shell_io_host_ar_bits_addr; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_r_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_host_r_valid; // @[DCRAccel.scala 53:21]
  wire [63:0] shell_io_host_r_bits_data; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_aw_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_aw_valid; // @[DCRAccel.scala 53:21]
  wire [31:0] shell_io_mem_aw_bits_addr; // @[DCRAccel.scala 53:21]
  wire [31:0] shell_io_mem_aw_bits_len; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_w_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_w_valid; // @[DCRAccel.scala 53:21]
  wire [63:0] shell_io_mem_w_bits_data; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_w_bits_last; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_b_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_b_valid; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_ar_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_ar_valid; // @[DCRAccel.scala 53:21]
  wire [31:0] shell_io_mem_ar_bits_addr; // @[DCRAccel.scala 53:21]
  wire [31:0] shell_io_mem_ar_bits_len; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_r_ready; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_r_valid; // @[DCRAccel.scala 53:21]
  wire [63:0] shell_io_mem_r_bits_data; // @[DCRAccel.scala 53:21]
  wire  shell_io_mem_r_bits_last; // @[DCRAccel.scala 53:21]
  AXISimShell sim_shell ( // @[DCRAccel.scala 52:25]
    .clock(sim_shell_clock),
    .reset(sim_shell_reset),
    .mem_aw_ready(sim_shell_mem_aw_ready),
    .mem_aw_valid(sim_shell_mem_aw_valid),
    .mem_aw_bits_addr(sim_shell_mem_aw_bits_addr),
    .mem_aw_bits_len(sim_shell_mem_aw_bits_len),
    .mem_w_ready(sim_shell_mem_w_ready),
    .mem_w_valid(sim_shell_mem_w_valid),
    .mem_w_bits_data(sim_shell_mem_w_bits_data),
    .mem_w_bits_last(sim_shell_mem_w_bits_last),
    .mem_b_ready(sim_shell_mem_b_ready),
    .mem_b_valid(sim_shell_mem_b_valid),
    .mem_ar_ready(sim_shell_mem_ar_ready),
    .mem_ar_valid(sim_shell_mem_ar_valid),
    .mem_ar_bits_addr(sim_shell_mem_ar_bits_addr),
    .mem_ar_bits_len(sim_shell_mem_ar_bits_len),
    .mem_r_ready(sim_shell_mem_r_ready),
    .mem_r_valid(sim_shell_mem_r_valid),
    .mem_r_bits_data(sim_shell_mem_r_bits_data),
    .mem_r_bits_last(sim_shell_mem_r_bits_last),
    .host_aw_ready(sim_shell_host_aw_ready),
    .host_aw_valid(sim_shell_host_aw_valid),
    .host_aw_bits_addr(sim_shell_host_aw_bits_addr),
    .host_w_ready(sim_shell_host_w_ready),
    .host_w_valid(sim_shell_host_w_valid),
    .host_w_bits_data(sim_shell_host_w_bits_data),
    .host_b_ready(sim_shell_host_b_ready),
    .host_b_valid(sim_shell_host_b_valid),
    .host_ar_ready(sim_shell_host_ar_ready),
    .host_ar_valid(sim_shell_host_ar_valid),
    .host_ar_bits_addr(sim_shell_host_ar_bits_addr),
    .host_r_ready(sim_shell_host_r_ready),
    .host_r_valid(sim_shell_host_r_valid),
    .host_r_bits_data(sim_shell_host_r_bits_data),
    .sim_clock(sim_shell_sim_clock),
    .sim_wait(sim_shell_sim_wait)
  );
  memGenDCRCacheShell shell ( // @[DCRAccel.scala 53:21]
    .clock(shell_clock),
    .reset(shell_reset),
    .io_host_aw_ready(shell_io_host_aw_ready),
    .io_host_aw_valid(shell_io_host_aw_valid),
    .io_host_aw_bits_addr(shell_io_host_aw_bits_addr),
    .io_host_w_ready(shell_io_host_w_ready),
    .io_host_w_valid(shell_io_host_w_valid),
    .io_host_w_bits_data(shell_io_host_w_bits_data),
    .io_host_b_ready(shell_io_host_b_ready),
    .io_host_b_valid(shell_io_host_b_valid),
    .io_host_ar_ready(shell_io_host_ar_ready),
    .io_host_ar_valid(shell_io_host_ar_valid),
    .io_host_ar_bits_addr(shell_io_host_ar_bits_addr),
    .io_host_r_ready(shell_io_host_r_ready),
    .io_host_r_valid(shell_io_host_r_valid),
    .io_host_r_bits_data(shell_io_host_r_bits_data),
    .io_mem_aw_ready(shell_io_mem_aw_ready),
    .io_mem_aw_valid(shell_io_mem_aw_valid),
    .io_mem_aw_bits_addr(shell_io_mem_aw_bits_addr),
    .io_mem_aw_bits_len(shell_io_mem_aw_bits_len),
    .io_mem_w_ready(shell_io_mem_w_ready),
    .io_mem_w_valid(shell_io_mem_w_valid),
    .io_mem_w_bits_data(shell_io_mem_w_bits_data),
    .io_mem_w_bits_last(shell_io_mem_w_bits_last),
    .io_mem_b_ready(shell_io_mem_b_ready),
    .io_mem_b_valid(shell_io_mem_b_valid),
    .io_mem_ar_ready(shell_io_mem_ar_ready),
    .io_mem_ar_valid(shell_io_mem_ar_valid),
    .io_mem_ar_bits_addr(shell_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(shell_io_mem_ar_bits_len),
    .io_mem_r_ready(shell_io_mem_r_ready),
    .io_mem_r_valid(shell_io_mem_r_valid),
    .io_mem_r_bits_data(shell_io_mem_r_bits_data),
    .io_mem_r_bits_last(shell_io_mem_r_bits_last)
  );
  assign sim_wait = sim_shell_sim_wait; // @[DCRAccel.scala 56:12]
  assign sim_shell_clock = clock;
  assign sim_shell_reset = reset;
  assign sim_shell_mem_aw_valid = shell_io_mem_aw_valid; // @[DCRAccel.scala 62:20]
  assign sim_shell_mem_aw_bits_addr = shell_io_mem_aw_bits_addr; // @[DCRAccel.scala 62:20]
  assign sim_shell_mem_aw_bits_len = shell_io_mem_aw_bits_len; // @[DCRAccel.scala 62:20]
  assign sim_shell_mem_w_valid = shell_io_mem_w_valid; // @[DCRAccel.scala 63:19]
  assign sim_shell_mem_w_bits_data = shell_io_mem_w_bits_data; // @[DCRAccel.scala 63:19]
  assign sim_shell_mem_w_bits_last = shell_io_mem_w_bits_last; // @[DCRAccel.scala 63:19]
  assign sim_shell_mem_b_ready = shell_io_mem_b_ready; // @[DCRAccel.scala 64:18]
  assign sim_shell_mem_ar_valid = shell_io_mem_ar_valid; // @[DCRAccel.scala 61:20]
  assign sim_shell_mem_ar_bits_addr = shell_io_mem_ar_bits_addr; // @[DCRAccel.scala 61:20]
  assign sim_shell_mem_ar_bits_len = shell_io_mem_ar_bits_len; // @[DCRAccel.scala 61:20]
  assign sim_shell_mem_r_ready = shell_io_mem_r_ready; // @[DCRAccel.scala 65:18]
  assign sim_shell_host_aw_ready = shell_io_host_aw_ready; // @[DCRAccel.scala 70:20]
  assign sim_shell_host_w_ready = shell_io_host_w_ready; // @[DCRAccel.scala 71:19]
  assign sim_shell_host_b_valid = shell_io_host_b_valid; // @[DCRAccel.scala 67:20]
  assign sim_shell_host_ar_ready = shell_io_host_ar_ready; // @[DCRAccel.scala 69:20]
  assign sim_shell_host_r_valid = shell_io_host_r_valid; // @[DCRAccel.scala 68:20]
  assign sim_shell_host_r_bits_data = shell_io_host_r_bits_data; // @[DCRAccel.scala 68:20]
  assign sim_shell_sim_clock = sim_clock; // @[DCRAccel.scala 55:23]
  assign shell_clock = clock;
  assign shell_reset = reset;
  assign shell_io_host_aw_valid = sim_shell_host_aw_valid; // @[DCRAccel.scala 70:20]
  assign shell_io_host_aw_bits_addr = sim_shell_host_aw_bits_addr; // @[DCRAccel.scala 70:20]
  assign shell_io_host_w_valid = sim_shell_host_w_valid; // @[DCRAccel.scala 71:19]
  assign shell_io_host_w_bits_data = sim_shell_host_w_bits_data; // @[DCRAccel.scala 71:19]
  assign shell_io_host_b_ready = sim_shell_host_b_ready; // @[DCRAccel.scala 67:20]
  assign shell_io_host_ar_valid = sim_shell_host_ar_valid; // @[DCRAccel.scala 69:20]
  assign shell_io_host_ar_bits_addr = sim_shell_host_ar_bits_addr; // @[DCRAccel.scala 69:20]
  assign shell_io_host_r_ready = sim_shell_host_r_ready; // @[DCRAccel.scala 68:20]
  assign shell_io_mem_aw_ready = sim_shell_mem_aw_ready; // @[DCRAccel.scala 62:20]
  assign shell_io_mem_w_ready = sim_shell_mem_w_ready; // @[DCRAccel.scala 63:19]
  assign shell_io_mem_b_valid = sim_shell_mem_b_valid; // @[DCRAccel.scala 64:18]
  assign shell_io_mem_ar_ready = sim_shell_mem_ar_ready; // @[DCRAccel.scala 61:20]
  assign shell_io_mem_r_valid = sim_shell_mem_r_valid; // @[DCRAccel.scala 65:18]
  assign shell_io_mem_r_bits_data = sim_shell_mem_r_bits_data; // @[DCRAccel.scala 65:18]
  assign shell_io_mem_r_bits_last = sim_shell_mem_r_bits_last; // @[DCRAccel.scala 65:18]
endmodule
